`timescale 1ns / 1fs 
module test_aes_128; 
reg clk; 
reg [127:0] state; 
reg [127:0] key; 
reg rst; 
wire [127:0] out; 
wire Antena; 
reg [127:0] bit_err; 
integer i; 
integer f; 
reg [127:0] out1; 
reg [127:0] out2; 
reg [127:0] out3; 
reg [127:0] out4; 
reg [127:0] out5; 
reg [127:0] out6; 
reg [127:0] out7; 
reg [127:0] out8; 
reg [127:0] out9; 
reg [127:0] out10; 
reg [127:0] out11; 
reg [127:0] out12; 
reg [127:0] out13; 
reg [127:0] out14; 
reg [127:0] out15; 
reg [127:0] out16; 
reg [127:0] out17; 
reg [127:0] out18; 
reg [127:0] out19; 
reg [127:0] out20; 
reg [127:0] out21; 
reg [127:0] out22; 
reg [127:0] out23; 
reg [127:0] out24; 
reg [127:0] out25; 
reg [127:0] out26; 
reg [127:0] out27; 
reg [127:0] out28; 
reg [127:0] out29; 
reg [127:0] out30; 
reg [127:0] out31; 
reg [127:0] out32; 
reg [127:0] out33; 
reg [127:0] out34; 
reg [127:0] out35; 
reg [127:0] out36; 
reg [127:0] out37; 
reg [127:0] out38; 
reg [127:0] out39; 
reg [127:0] out40; 
reg [127:0] out41; 
reg [127:0] out42; 
reg [127:0] out43; 
reg [127:0] out44; 
reg [127:0] out45; 
reg [127:0] out46; 
reg [127:0] out47; 
reg [127:0] out48; 
reg [127:0] out49; 
reg [127:0] out50; 
reg [127:0] out51; 
reg [127:0] out52; 
reg [127:0] out53; 
reg [127:0] out54; 
reg [127:0] out55; 
reg [127:0] out56; 
reg [127:0] out57; 
reg [127:0] out58; 
reg [127:0] out59; 
reg [127:0] out60; 
reg [127:0] out61; 
reg [127:0] out62; 
reg [127:0] out63; 
reg [127:0] out64; 
reg [127:0] out65; 
reg [127:0] out66; 
reg [127:0] out67; 
reg [127:0] out68; 
reg [127:0] out69; 
reg [127:0] out70; 
reg [127:0] out71; 
reg [127:0] out72; 
reg [127:0] out73; 
reg [127:0] out74; 
reg [127:0] out75; 
reg [127:0] out76; 
reg [127:0] out77; 
reg [127:0] out78; 
reg [127:0] out79; 
reg [127:0] out80; 
reg [127:0] out81; 
reg [127:0] out82; 
reg [127:0] out83; 
reg [127:0] out84; 
reg [127:0] out85; 
reg [127:0] out86; 
reg [127:0] out87; 
reg [127:0] out88; 
reg [127:0] out89; 
reg [127:0] out90; 
reg [127:0] out91; 
reg [127:0] out92; 
reg [127:0] out93; 
reg [127:0] out94; 
reg [127:0] out95; 
reg [127:0] out96; 
reg [127:0] out97; 
reg [127:0] out98; 
reg [127:0] out99; 
reg [127:0] out100; 
reg [127:0] out101; 
reg [127:0] out102; 
reg [127:0] out103; 
reg [127:0] out104; 
reg [127:0] out105; 
reg [127:0] out106; 
reg [127:0] out107; 
reg [127:0] out108; 
reg [127:0] out109; 
reg [127:0] out110; 
reg [127:0] out111; 
reg [127:0] out112; 
reg [127:0] out113; 
reg [127:0] out114; 
reg [127:0] out115; 
reg [127:0] out116; 
reg [127:0] out117; 
reg [127:0] out118; 
reg [127:0] out119; 
reg [127:0] out120; 
reg [127:0] out121; 
reg [127:0] out122; 
reg [127:0] out123; 
reg [127:0] out124; 
reg [127:0] out125; 
reg [127:0] out126; 
reg [127:0] out127; 
reg [127:0] out128; 
reg [127:0] out129; 
reg [127:0] out130; 
reg [127:0] out131; 
reg [127:0] out132; 
reg [127:0] out133; 
reg [127:0] out134; 
reg [127:0] out135; 
reg [127:0] out136; 
reg [127:0] out137; 
reg [127:0] out138; 
reg [127:0] out139; 
reg [127:0] out140; 
reg [127:0] out141; 
reg [127:0] out142; 
reg [127:0] out143; 
reg [127:0] out144; 
reg [127:0] out145; 
reg [127:0] out146; 
reg [127:0] out147; 
reg [127:0] out148; 
reg [127:0] out149; 
reg [127:0] out150; 
reg [127:0] out151; 
reg [127:0] out152; 
reg [127:0] out153; 
reg [127:0] out154; 
reg [127:0] out155; 
reg [127:0] out156; 
reg [127:0] out157; 
reg [127:0] out158; 
reg [127:0] out159; 
reg [127:0] out160; 
reg [127:0] out161; 
reg [127:0] out162; 
reg [127:0] out163; 
reg [127:0] out164; 
reg [127:0] out165; 
reg [127:0] out166; 
reg [127:0] out167; 
reg [127:0] out168; 
reg [127:0] out169; 
reg [127:0] out170; 
reg [127:0] out171; 
reg [127:0] out172; 
reg [127:0] out173; 
reg [127:0] out174; 
reg [127:0] out175; 
reg [127:0] out176; 
reg [127:0] out177; 
reg [127:0] out178; 
reg [127:0] out179; 
reg [127:0] out180; 
reg [127:0] out181; 
reg [127:0] out182; 
reg [127:0] out183; 
reg [127:0] out184; 
reg [127:0] out185; 
reg [127:0] out186; 
reg [127:0] out187; 
reg [127:0] out188; 
reg [127:0] out189; 
reg [127:0] out190; 
reg [127:0] out191; 
reg [127:0] out192; 
reg [127:0] out193; 
reg [127:0] out194; 
reg [127:0] out195; 
reg [127:0] out196; 
reg [127:0] out197; 
reg [127:0] out198; 
reg [127:0] out199; 
reg [127:0] out200; 
reg [127:0] out201; 
reg [127:0] out202; 
reg [127:0] out203; 
reg [127:0] out204; 
reg [127:0] out205; 
reg [127:0] out206; 
reg [127:0] out207; 
reg [127:0] out208; 
reg [127:0] out209; 
reg [127:0] out210; 
reg [127:0] out211; 
reg [127:0] out212; 
reg [127:0] out213; 
reg [127:0] out214; 
reg [127:0] out215; 
reg [127:0] out216; 
reg [127:0] out217; 
reg [127:0] out218; 
reg [127:0] out219; 
reg [127:0] out220; 
reg [127:0] out221; 
reg [127:0] out222; 
reg [127:0] out223; 
reg [127:0] out224; 
reg [127:0] out225; 
reg [127:0] out226; 
reg [127:0] out227; 
reg [127:0] out228; 
reg [127:0] out229; 
reg [127:0] out230; 
reg [127:0] out231; 
reg [127:0] out232; 
reg [127:0] out233; 
reg [127:0] out234; 
reg [127:0] out235; 
reg [127:0] out236; 
reg [127:0] out237; 
reg [127:0] out238; 
reg [127:0] out239; 
reg [127:0] out240; 
reg [127:0] out241; 
reg [127:0] out242; 
reg [127:0] out243; 
reg [127:0] out244; 
reg [127:0] out245; 
reg [127:0] out246; 
reg [127:0] out247; 
reg [127:0] out248; 
reg [127:0] out249; 
reg [127:0] out250; 
reg [127:0] out251; 
reg [127:0] out252; 
reg [127:0] out253; 
reg [127:0] out254; 
reg [127:0] out255; 
reg [127:0] out256; 
reg [127:0] out257; 
reg [127:0] out258; 
reg [127:0] out259; 
reg [127:0] out260; 
reg [127:0] out261; 
reg [127:0] out262; 
reg [127:0] out263; 
reg [127:0] out264; 
reg [127:0] out265; 
reg [127:0] out266; 
reg [127:0] out267; 
reg [127:0] out268; 
reg [127:0] out269; 
reg [127:0] out270; 
reg [127:0] out271; 
reg [127:0] out272; 
reg [127:0] out273; 
reg [127:0] out274; 
reg [127:0] out275; 
reg [127:0] out276; 
reg [127:0] out277; 
reg [127:0] out278; 
reg [127:0] out279; 
reg [127:0] out280; 
reg [127:0] out281; 
reg [127:0] out282; 
reg [127:0] out283; 
reg [127:0] out284; 
reg [127:0] out285; 
reg [127:0] out286; 
reg [127:0] out287; 
reg [127:0] out288; 
reg [127:0] out289; 
reg [127:0] out290; 
reg [127:0] out291; 
reg [127:0] out292; 
reg [127:0] out293; 
reg [127:0] out294; 
reg [127:0] out295; 
reg [127:0] out296; 
reg [127:0] out297; 
reg [127:0] out298; 
reg [127:0] out299; 
reg [127:0] out300; 
reg [127:0] out301; 
reg [127:0] out302; 
reg [127:0] out303; 
reg [127:0] out304; 
reg [127:0] out305; 
reg [127:0] out306; 
reg [127:0] out307; 
reg [127:0] out308; 
reg [127:0] out309; 
reg [127:0] out310; 
reg [127:0] out311; 
reg [127:0] out312; 
reg [127:0] out313; 
reg [127:0] out314; 
reg [127:0] out315; 
reg [127:0] out316; 
reg [127:0] out317; 
reg [127:0] out318; 
reg [127:0] out319; 
reg [127:0] out320; 
reg [127:0] out321; 
reg [127:0] out322; 
reg [127:0] out323; 
reg [127:0] out324; 
reg [127:0] out325; 
reg [127:0] out326; 
reg [127:0] out327; 
reg [127:0] out328; 
reg [127:0] out329; 
reg [127:0] out330; 
reg [127:0] out331; 
reg [127:0] out332; 
reg [127:0] out333; 
reg [127:0] out334; 
reg [127:0] out335; 
reg [127:0] out336; 
reg [127:0] out337; 
reg [127:0] out338; 
reg [127:0] out339; 
reg [127:0] out340; 
reg [127:0] out341; 
reg [127:0] out342; 
reg [127:0] out343; 
reg [127:0] out344; 
reg [127:0] out345; 
reg [127:0] out346; 
reg [127:0] out347; 
reg [127:0] out348; 
reg [127:0] out349; 
reg [127:0] out350; 
reg [127:0] out351; 
reg [127:0] out352; 
reg [127:0] out353; 
reg [127:0] out354; 
reg [127:0] out355; 
reg [127:0] out356; 
reg [127:0] out357; 
reg [127:0] out358; 
reg [127:0] out359; 
reg [127:0] out360; 
reg [127:0] out361; 
reg [127:0] out362; 
reg [127:0] out363; 
reg [127:0] out364; 
reg [127:0] out365; 
reg [127:0] out366; 
reg [127:0] out367; 
reg [127:0] out368; 
reg [127:0] out369; 
reg [127:0] out370; 
reg [127:0] out371; 
reg [127:0] out372; 
reg [127:0] out373; 
reg [127:0] out374; 
reg [127:0] out375; 
reg [127:0] out376; 
reg [127:0] out377; 
reg [127:0] out378; 
reg [127:0] out379; 
reg [127:0] out380; 
reg [127:0] out381; 
reg [127:0] out382; 
reg [127:0] out383; 
reg [127:0] out384; 
reg [127:0] out385; 
reg [127:0] out386; 
reg [127:0] out387; 
reg [127:0] out388; 
reg [127:0] out389; 
reg [127:0] out390; 
reg [127:0] out391; 
reg [127:0] out392; 
reg [127:0] out393; 
reg [127:0] out394; 
reg [127:0] out395; 
reg [127:0] out396; 
reg [127:0] out397; 
reg [127:0] out398; 
reg [127:0] out399; 
reg [127:0] out400; 
reg [127:0] out401; 
reg [127:0] out402; 
reg [127:0] out403; 
reg [127:0] out404; 
reg [127:0] out405; 
reg [127:0] out406; 
reg [127:0] out407; 
reg [127:0] out408; 
reg [127:0] out409; 
reg [127:0] out410; 
reg [127:0] out411; 
reg [127:0] out412; 
reg [127:0] out413; 
reg [127:0] out414; 
reg [127:0] out415; 
reg [127:0] out416; 
reg [127:0] out417; 
reg [127:0] out418; 
reg [127:0] out419; 
reg [127:0] out420; 
reg [127:0] out421; 
reg [127:0] out422; 
reg [127:0] out423; 
reg [127:0] out424; 
reg [127:0] out425; 
reg [127:0] out426; 
reg [127:0] out427; 
reg [127:0] out428; 
reg [127:0] out429; 
reg [127:0] out430; 
reg [127:0] out431; 
reg [127:0] out432; 
reg [127:0] out433; 
reg [127:0] out434; 
reg [127:0] out435; 
reg [127:0] out436; 
reg [127:0] out437; 
reg [127:0] out438; 
reg [127:0] out439; 
reg [127:0] out440; 
reg [127:0] out441; 
reg [127:0] out442; 
reg [127:0] out443; 
reg [127:0] out444; 
reg [127:0] out445; 
reg [127:0] out446; 
reg [127:0] out447; 
reg [127:0] out448; 
reg [127:0] out449; 
reg [127:0] out450; 
reg [127:0] out451; 
reg [127:0] out452; 
reg [127:0] out453; 
reg [127:0] out454; 
reg [127:0] out455; 
reg [127:0] out456; 
reg [127:0] out457; 
reg [127:0] out458; 
reg [127:0] out459; 
reg [127:0] out460; 
reg [127:0] out461; 
reg [127:0] out462; 
reg [127:0] out463; 
reg [127:0] out464; 
reg [127:0] out465; 
reg [127:0] out466; 
reg [127:0] out467; 
reg [127:0] out468; 
reg [127:0] out469; 
reg [127:0] out470; 
reg [127:0] out471; 
reg [127:0] out472; 
reg [127:0] out473; 
reg [127:0] out474; 
reg [127:0] out475; 
reg [127:0] out476; 
reg [127:0] out477; 
reg [127:0] out478; 
reg [127:0] out479; 
reg [127:0] out480; 
reg [127:0] out481; 
reg [127:0] out482; 
reg [127:0] out483; 
reg [127:0] out484; 
reg [127:0] out485; 
reg [127:0] out486; 
reg [127:0] out487; 
reg [127:0] out488; 
reg [127:0] out489; 
reg [127:0] out490; 
reg [127:0] out491; 
reg [127:0] out492; 
reg [127:0] out493; 
reg [127:0] out494; 
reg [127:0] out495; 
reg [127:0] out496; 
reg [127:0] out497; 
reg [127:0] out498; 
reg [127:0] out499; 
reg [127:0] out500; 
reg [127:0] out501; 
reg [127:0] out502; 
reg [127:0] out503; 
reg [127:0] out504; 
reg [127:0] out505; 
reg [127:0] out506; 
reg [127:0] out507; 
reg [127:0] out508; 
reg [127:0] out509; 
reg [127:0] out510; 
reg [127:0] out511; 
reg [127:0] out512; 
reg [127:0] out513; 
reg [127:0] out514; 
reg [127:0] out515; 
reg [127:0] out516; 
reg [127:0] out517; 
reg [127:0] out518; 
reg [127:0] out519; 
reg [127:0] out520; 
reg [127:0] out521; 
reg [127:0] out522; 
reg [127:0] out523; 
reg [127:0] out524; 
reg [127:0] out525; 
reg [127:0] out526; 
reg [127:0] out527; 
reg [127:0] out528; 
reg [127:0] out529; 
reg [127:0] out530; 
reg [127:0] out531; 
reg [127:0] out532; 
reg [127:0] out533; 
reg [127:0] out534; 
reg [127:0] out535; 
reg [127:0] out536; 
reg [127:0] out537; 
reg [127:0] out538; 
reg [127:0] out539; 
reg [127:0] out540; 
reg [127:0] out541; 
reg [127:0] out542; 
reg [127:0] out543; 
reg [127:0] out544; 
reg [127:0] out545; 
reg [127:0] out546; 
reg [127:0] out547; 
reg [127:0] out548; 
reg [127:0] out549; 
reg [127:0] out550; 
reg [127:0] out551; 
reg [127:0] out552; 
reg [127:0] out553; 
reg [127:0] out554; 
reg [127:0] out555; 
reg [127:0] out556; 
reg [127:0] out557; 
reg [127:0] out558; 
reg [127:0] out559; 
reg [127:0] out560; 
reg [127:0] out561; 
reg [127:0] out562; 
reg [127:0] out563; 
reg [127:0] out564; 
reg [127:0] out565; 
reg [127:0] out566; 
reg [127:0] out567; 
reg [127:0] out568; 
reg [127:0] out569; 
reg [127:0] out570; 
reg [127:0] out571; 
reg [127:0] out572; 
reg [127:0] out573; 
reg [127:0] out574; 
reg [127:0] out575; 
reg [127:0] out576; 
reg [127:0] out577; 
reg [127:0] out578; 
reg [127:0] out579; 
reg [127:0] out580; 
reg [127:0] out581; 
reg [127:0] out582; 
reg [127:0] out583; 
reg [127:0] out584; 
reg [127:0] out585; 
reg [127:0] out586; 
reg [127:0] out587; 
reg [127:0] out588; 
reg [127:0] out589; 
reg [127:0] out590; 
reg [127:0] out591; 
reg [127:0] out592; 
reg [127:0] out593; 
reg [127:0] out594; 
reg [127:0] out595; 
reg [127:0] out596; 
reg [127:0] out597; 
reg [127:0] out598; 
reg [127:0] out599; 
reg [127:0] out600; 
reg [127:0] out601; 
reg [127:0] out602; 
reg [127:0] out603; 
reg [127:0] out604; 
reg [127:0] out605; 
reg [127:0] out606; 
reg [127:0] out607; 
reg [127:0] out608; 
reg [127:0] out609; 
reg [127:0] out610; 
reg [127:0] out611; 
reg [127:0] out612; 
reg [127:0] out613; 
reg [127:0] out614; 
reg [127:0] out615; 
reg [127:0] out616; 
reg [127:0] out617; 
reg [127:0] out618; 
reg [127:0] out619; 
reg [127:0] out620; 
reg [127:0] out621; 
reg [127:0] out622; 
reg [127:0] out623; 
reg [127:0] out624; 
reg [127:0] out625; 
reg [127:0] out626; 
reg [127:0] out627; 
reg [127:0] out628; 
reg [127:0] out629; 
reg [127:0] out630; 
reg [127:0] out631; 
reg [127:0] out632; 
reg [127:0] out633; 
reg [127:0] out634; 
reg [127:0] out635; 
reg [127:0] out636; 
reg [127:0] out637; 
reg [127:0] out638; 
reg [127:0] out639; 
reg [127:0] out640; 
reg [127:0] out641; 
reg [127:0] out642; 
reg [127:0] out643; 
reg [127:0] out644; 
reg [127:0] out645; 
reg [127:0] out646; 
reg [127:0] out647; 
reg [127:0] out648; 
reg [127:0] out649; 
reg [127:0] out650; 
reg [127:0] out651; 
reg [127:0] out652; 
reg [127:0] out653; 
reg [127:0] out654; 
reg [127:0] out655; 
reg [127:0] out656; 
reg [127:0] out657; 
reg [127:0] out658; 
reg [127:0] out659; 
reg [127:0] out660; 
reg [127:0] out661; 
reg [127:0] out662; 
reg [127:0] out663; 
reg [127:0] out664; 
reg [127:0] out665; 
reg [127:0] out666; 
reg [127:0] out667; 
reg [127:0] out668; 
reg [127:0] out669; 
reg [127:0] out670; 
reg [127:0] out671; 
reg [127:0] out672; 
reg [127:0] out673; 
reg [127:0] out674; 
reg [127:0] out675; 
reg [127:0] out676; 
reg [127:0] out677; 
reg [127:0] out678; 
reg [127:0] out679; 
reg [127:0] out680; 
reg [127:0] out681; 
reg [127:0] out682; 
reg [127:0] out683; 
reg [127:0] out684; 
reg [127:0] out685; 
reg [127:0] out686; 
reg [127:0] out687; 
reg [127:0] out688; 
reg [127:0] out689; 
reg [127:0] out690; 
reg [127:0] out691; 
reg [127:0] out692; 
reg [127:0] out693; 
reg [127:0] out694; 
reg [127:0] out695; 
reg [127:0] out696; 
reg [127:0] out697; 
reg [127:0] out698; 
reg [127:0] out699; 
reg [127:0] out700; 
reg [127:0] out701; 
reg [127:0] out702; 
reg [127:0] out703; 
reg [127:0] out704; 
reg [127:0] out705; 
reg [127:0] out706; 
reg [127:0] out707; 
reg [127:0] out708; 
reg [127:0] out709; 
reg [127:0] out710; 
reg [127:0] out711; 
reg [127:0] out712; 
reg [127:0] out713; 
reg [127:0] out714; 
reg [127:0] out715; 
reg [127:0] out716; 
reg [127:0] out717; 
reg [127:0] out718; 
reg [127:0] out719; 
reg [127:0] out720; 
reg [127:0] out721; 
reg [127:0] out722; 
reg [127:0] out723; 
reg [127:0] out724; 
reg [127:0] out725; 
reg [127:0] out726; 
reg [127:0] out727; 
reg [127:0] out728; 
reg [127:0] out729; 
reg [127:0] out730; 
reg [127:0] out731; 
reg [127:0] out732; 
reg [127:0] out733; 
reg [127:0] out734; 
reg [127:0] out735; 
reg [127:0] out736; 
reg [127:0] out737; 
reg [127:0] out738; 
reg [127:0] out739; 
reg [127:0] out740; 
reg [127:0] out741; 
reg [127:0] out742; 
reg [127:0] out743; 
reg [127:0] out744; 
reg [127:0] out745; 
reg [127:0] out746; 
reg [127:0] out747; 
reg [127:0] out748; 
reg [127:0] out749; 
reg [127:0] out750; 
reg [127:0] out751; 
reg [127:0] out752; 
reg [127:0] out753; 
reg [127:0] out754; 
reg [127:0] out755; 
reg [127:0] out756; 
reg [127:0] out757; 
reg [127:0] out758; 
reg [127:0] out759; 
reg [127:0] out760; 
reg [127:0] out761; 
reg [127:0] out762; 
reg [127:0] out763; 
reg [127:0] out764; 
reg [127:0] out765; 
reg [127:0] out766; 
reg [127:0] out767; 
reg [127:0] out768; 
reg [127:0] out769; 
reg [127:0] out770; 
reg [127:0] out771; 
reg [127:0] out772; 
reg [127:0] out773; 
reg [127:0] out774; 
reg [127:0] out775; 
reg [127:0] out776; 
reg [127:0] out777; 
reg [127:0] out778; 
reg [127:0] out779; 
reg [127:0] out780; 
reg [127:0] out781; 
reg [127:0] out782; 
reg [127:0] out783; 
reg [127:0] out784; 
reg [127:0] out785; 
reg [127:0] out786; 
reg [127:0] out787; 
reg [127:0] out788; 
reg [127:0] out789; 
reg [127:0] out790; 
reg [127:0] out791; 
reg [127:0] out792; 
reg [127:0] out793; 
reg [127:0] out794; 
reg [127:0] out795; 
reg [127:0] out796; 
reg [127:0] out797; 
reg [127:0] out798; 
reg [127:0] out799; 
reg [127:0] out800; 
reg [127:0] out801; 
reg [127:0] out802; 
reg [127:0] out803; 
reg [127:0] out804; 
reg [127:0] out805; 
reg [127:0] out806; 
reg [127:0] out807; 
reg [127:0] out808; 
reg [127:0] out809; 
reg [127:0] out810; 
reg [127:0] out811; 
reg [127:0] out812; 
reg [127:0] out813; 
reg [127:0] out814; 
reg [127:0] out815; 
reg [127:0] out816; 
reg [127:0] out817; 
reg [127:0] out818; 
reg [127:0] out819; 
reg [127:0] out820; 
reg [127:0] out821; 
reg [127:0] out822; 
reg [127:0] out823; 
reg [127:0] out824; 
reg [127:0] out825; 
reg [127:0] out826; 
reg [127:0] out827; 
reg [127:0] out828; 
reg [127:0] out829; 
reg [127:0] out830; 
reg [127:0] out831; 
reg [127:0] out832; 
reg [127:0] out833; 
reg [127:0] out834; 
reg [127:0] out835; 
reg [127:0] out836; 
reg [127:0] out837; 
reg [127:0] out838; 
reg [127:0] out839; 
reg [127:0] out840; 
reg [127:0] out841; 
reg [127:0] out842; 
reg [127:0] out843; 
reg [127:0] out844; 
reg [127:0] out845; 
reg [127:0] out846; 
reg [127:0] out847; 
reg [127:0] out848; 
reg [127:0] out849; 
reg [127:0] out850; 
reg [127:0] out851; 
reg [127:0] out852; 
reg [127:0] out853; 
reg [127:0] out854; 
reg [127:0] out855; 
reg [127:0] out856; 
reg [127:0] out857; 
reg [127:0] out858; 
reg [127:0] out859; 
reg [127:0] out860; 
reg [127:0] out861; 
reg [127:0] out862; 
reg [127:0] out863; 
reg [127:0] out864; 
reg [127:0] out865; 
reg [127:0] out866; 
reg [127:0] out867; 
reg [127:0] out868; 
reg [127:0] out869; 
reg [127:0] out870; 
reg [127:0] out871; 
reg [127:0] out872; 
reg [127:0] out873; 
reg [127:0] out874; 
reg [127:0] out875; 
reg [127:0] out876; 
reg [127:0] out877; 
reg [127:0] out878; 
reg [127:0] out879; 
reg [127:0] out880; 
reg [127:0] out881; 
reg [127:0] out882; 
reg [127:0] out883; 
reg [127:0] out884; 
reg [127:0] out885; 
reg [127:0] out886; 
reg [127:0] out887; 
reg [127:0] out888; 
reg [127:0] out889; 
reg [127:0] out890; 
reg [127:0] out891; 
reg [127:0] out892; 
reg [127:0] out893; 
reg [127:0] out894; 
reg [127:0] out895; 
reg [127:0] out896; 
reg [127:0] out897; 
reg [127:0] out898; 
reg [127:0] out899; 
reg [127:0] out900; 
reg [127:0] out901; 
reg [127:0] out902; 
reg [127:0] out903; 
reg [127:0] out904; 
reg [127:0] out905; 
reg [127:0] out906; 
reg [127:0] out907; 
reg [127:0] out908; 
reg [127:0] out909; 
reg [127:0] out910; 
reg [127:0] out911; 
reg [127:0] out912; 
reg [127:0] out913; 
reg [127:0] out914; 
reg [127:0] out915; 
reg [127:0] out916; 
reg [127:0] out917; 
reg [127:0] out918; 
reg [127:0] out919; 
reg [127:0] out920; 
reg [127:0] out921; 
reg [127:0] out922; 
reg [127:0] out923; 
reg [127:0] out924; 
reg [127:0] out925; 
reg [127:0] out926; 
reg [127:0] out927; 
reg [127:0] out928; 
reg [127:0] out929; 
reg [127:0] out930; 
reg [127:0] out931; 
reg [127:0] out932; 
reg [127:0] out933; 
reg [127:0] out934; 
reg [127:0] out935; 
reg [127:0] out936; 
reg [127:0] out937; 
reg [127:0] out938; 
reg [127:0] out939; 
reg [127:0] out940; 
reg [127:0] out941; 
reg [127:0] out942; 
reg [127:0] out943; 
reg [127:0] out944; 
reg [127:0] out945; 
reg [127:0] out946; 
reg [127:0] out947; 
reg [127:0] out948; 
reg [127:0] out949; 
reg [127:0] out950; 
reg [127:0] out951; 
reg [127:0] out952; 
reg [127:0] out953; 
reg [127:0] out954; 
reg [127:0] out955; 
reg [127:0] out956; 
reg [127:0] out957; 
reg [127:0] out958; 
reg [127:0] out959; 
reg [127:0] out960; 
reg [127:0] out961; 
reg [127:0] out962; 
reg [127:0] out963; 
reg [127:0] out964; 
reg [127:0] out965; 
reg [127:0] out966; 
reg [127:0] out967; 
reg [127:0] out968; 
reg [127:0] out969; 
reg [127:0] out970; 
reg [127:0] out971; 
reg [127:0] out972; 
reg [127:0] out973; 
reg [127:0] out974; 
reg [127:0] out975; 
reg [127:0] out976; 
reg [127:0] out977; 
reg [127:0] out978; 
reg [127:0] out979; 
reg [127:0] out980; 
reg [127:0] out981; 
reg [127:0] out982; 
reg [127:0] out983; 
reg [127:0] out984; 
reg [127:0] out985; 
reg [127:0] out986; 
reg [127:0] out987; 
reg [127:0] out988; 
reg [127:0] out989; 
reg [127:0] out990; 
reg [127:0] out991; 
reg [127:0] out992; 
reg [127:0] out993; 
reg [127:0] out994; 
reg [127:0] out995; 
reg [127:0] out996; 
reg [127:0] out997; 
reg [127:0] out998; 
reg [127:0] out999; 
reg [127:0] out1000; 
reg [127:0] out1001; 
reg [127:0] out1002; 
reg [127:0] out1003; 
reg [127:0] out1004; 
reg [127:0] out1005; 
reg [127:0] out1006; 
reg [127:0] out1007; 
reg [127:0] out1008; 
reg [127:0] out1009; 
reg [127:0] out1010; 
reg [127:0] out1011; 
reg [127:0] out1012; 
reg [127:0] out1013; 
reg [127:0] out1014; 
reg [127:0] out1015; 
reg [127:0] out1016; 
reg [127:0] out1017; 
reg [127:0] out1018; 
reg [127:0] out1019; 
reg [127:0] out1020; 
reg [127:0] out1021; 
reg [127:0] out1022; 
reg [127:0] out1023; 
reg [127:0] out1024; 
reg [127:0] out1025; 
reg [127:0] out1026; 
reg [127:0] out1027; 
reg [127:0] out1028; 
reg [127:0] out1029; 
reg [127:0] out1030; 
reg [127:0] out1031; 
reg [127:0] out1032; 
reg [127:0] out1033; 
reg [127:0] out1034; 
reg [127:0] out1035; 
reg [127:0] out1036; 
reg [127:0] out1037; 
reg [127:0] out1038; 
reg [127:0] out1039; 
reg [127:0] out1040; 
reg [127:0] out1041; 
reg [127:0] out1042; 
reg [127:0] out1043; 
reg [127:0] out1044; 
reg [127:0] out1045; 
reg [127:0] out1046; 
reg [127:0] out1047; 
reg [127:0] out1048; 
reg [127:0] out1049; 
reg [127:0] out1050; 
reg [127:0] out1051; 
reg [127:0] out1052; 
reg [127:0] out1053; 
reg [127:0] out1054; 
reg [127:0] out1055; 
reg [127:0] out1056; 
reg [127:0] out1057; 
reg [127:0] out1058; 
reg [127:0] out1059; 
reg [127:0] out1060; 
reg [127:0] out1061; 
reg [127:0] out1062; 
reg [127:0] out1063; 
reg [127:0] out1064; 
reg [127:0] out1065; 
reg [127:0] out1066; 
reg [127:0] out1067; 
reg [127:0] out1068; 
reg [127:0] out1069; 
reg [127:0] out1070; 
reg [127:0] out1071; 
reg [127:0] out1072; 
reg [127:0] out1073; 
reg [127:0] out1074; 
reg [127:0] out1075; 
reg [127:0] out1076; 
reg [127:0] out1077; 
reg [127:0] out1078; 
reg [127:0] out1079; 
reg [127:0] out1080; 
reg [127:0] out1081; 
reg [127:0] out1082; 
reg [127:0] out1083; 
reg [127:0] out1084; 
reg [127:0] out1085; 
reg [127:0] out1086; 
reg [127:0] out1087; 
reg [127:0] out1088; 
reg [127:0] out1089; 
reg [127:0] out1090; 
reg [127:0] out1091; 
reg [127:0] out1092; 
reg [127:0] out1093; 
reg [127:0] out1094; 
reg [127:0] out1095; 
reg [127:0] out1096; 
reg [127:0] out1097; 
reg [127:0] out1098; 
reg [127:0] out1099; 
reg [127:0] out1100; 
reg [127:0] out1101; 
reg [127:0] out1102; 
reg [127:0] out1103; 
reg [127:0] out1104; 
reg [127:0] out1105; 
reg [127:0] out1106; 
reg [127:0] out1107; 
reg [127:0] out1108; 
reg [127:0] out1109; 
reg [127:0] out1110; 
reg [127:0] out1111; 
reg [127:0] out1112; 
reg [127:0] out1113; 
reg [127:0] out1114; 
reg [127:0] out1115; 
reg [127:0] out1116; 
reg [127:0] out1117; 
reg [127:0] out1118; 
reg [127:0] out1119; 
reg [127:0] out1120; 
reg [127:0] out1121; 
reg [127:0] out1122; 
reg [127:0] out1123; 
reg [127:0] out1124; 
reg [127:0] out1125; 
reg [127:0] out1126; 
reg [127:0] out1127; 
reg [127:0] out1128; 
reg [127:0] out1129; 
reg [127:0] out1130; 
reg [127:0] out1131; 
reg [127:0] out1132; 
reg [127:0] out1133; 
reg [127:0] out1134; 
reg [127:0] out1135; 
reg [127:0] out1136; 
reg [127:0] out1137; 
reg [127:0] out1138; 
reg [127:0] out1139; 
reg [127:0] out1140; 
reg [127:0] out1141; 
reg [127:0] out1142; 
reg [127:0] out1143; 
reg [127:0] out1144; 
reg [127:0] out1145; 
reg [127:0] out1146; 
reg [127:0] out1147; 
reg [127:0] out1148; 
reg [127:0] out1149; 
reg [127:0] out1150; 
reg [127:0] out1151; 
reg [127:0] out1152; 
reg [127:0] out1153; 
reg [127:0] out1154; 
reg [127:0] out1155; 
reg [127:0] out1156; 
reg [127:0] out1157; 
reg [127:0] out1158; 
reg [127:0] out1159; 
reg [127:0] out1160; 
reg [127:0] out1161; 
reg [127:0] out1162; 
reg [127:0] out1163; 
reg [127:0] out1164; 
reg [127:0] out1165; 
reg [127:0] out1166; 
reg [127:0] out1167; 
reg [127:0] out1168; 
reg [127:0] out1169; 
reg [127:0] out1170; 
reg [127:0] out1171; 
reg [127:0] out1172; 
reg [127:0] out1173; 
reg [127:0] out1174; 
reg [127:0] out1175; 
reg [127:0] out1176; 
reg [127:0] out1177; 
reg [127:0] out1178; 
reg [127:0] out1179; 
reg [127:0] out1180; 
reg [127:0] out1181; 
reg [127:0] out1182; 
reg [127:0] out1183; 
reg [127:0] out1184; 
reg [127:0] out1185; 
reg [127:0] out1186; 
reg [127:0] out1187; 
reg [127:0] out1188; 
reg [127:0] out1189; 
reg [127:0] out1190; 
reg [127:0] out1191; 
reg [127:0] out1192; 
reg [127:0] out1193; 
reg [127:0] out1194; 
reg [127:0] out1195; 
reg [127:0] out1196; 
reg [127:0] out1197; 
reg [127:0] out1198; 
reg [127:0] out1199; 
reg [127:0] out1200; 
reg [127:0] out1201; 
reg [127:0] out1202; 
reg [127:0] out1203; 
reg [127:0] out1204; 
reg [127:0] out1205; 
reg [127:0] out1206; 
reg [127:0] out1207; 
reg [127:0] out1208; 
reg [127:0] out1209; 
reg [127:0] out1210; 
reg [127:0] out1211; 
reg [127:0] out1212; 
reg [127:0] out1213; 
reg [127:0] out1214; 
reg [127:0] out1215; 
reg [127:0] out1216; 
reg [127:0] out1217; 
reg [127:0] out1218; 
reg [127:0] out1219; 
reg [127:0] out1220; 
reg [127:0] out1221; 
reg [127:0] out1222; 
reg [127:0] out1223; 
reg [127:0] out1224; 
reg [127:0] out1225; 
reg [127:0] out1226; 
reg [127:0] out1227; 
reg [127:0] out1228; 
reg [127:0] out1229; 
reg [127:0] out1230; 
reg [127:0] out1231; 
reg [127:0] out1232; 
reg [127:0] out1233; 
reg [127:0] out1234; 
reg [127:0] out1235; 
reg [127:0] out1236; 
reg [127:0] out1237; 
reg [127:0] out1238; 
reg [127:0] out1239; 
reg [127:0] out1240; 
reg [127:0] out1241; 
reg [127:0] out1242; 
reg [127:0] out1243; 
reg [127:0] out1244; 
reg [127:0] out1245; 
reg [127:0] out1246; 
reg [127:0] out1247; 
reg [127:0] out1248; 
reg [127:0] out1249; 
reg [127:0] out1250; 
reg [127:0] out1251; 
reg [127:0] out1252; 
reg [127:0] out1253; 
reg [127:0] out1254; 
reg [127:0] out1255; 
reg [127:0] out1256; 
reg [127:0] out1257; 
reg [127:0] out1258; 
reg [127:0] out1259; 
reg [127:0] out1260; 
reg [127:0] out1261; 
reg [127:0] out1262; 
reg [127:0] out1263; 
reg [127:0] out1264; 
reg [127:0] out1265; 
reg [127:0] out1266; 
reg [127:0] out1267; 
reg [127:0] out1268; 
reg [127:0] out1269; 
reg [127:0] out1270; 
reg [127:0] out1271; 
reg [127:0] out1272; 
reg [127:0] out1273; 
reg [127:0] out1274; 
reg [127:0] out1275; 
reg [127:0] out1276; 
reg [127:0] out1277; 
reg [127:0] out1278; 
reg [127:0] out1279; 
reg [127:0] out1280; 
reg [127:0] out1281; 
reg [127:0] out1282; 
reg [127:0] out1283; 
reg [127:0] out1284; 
reg [127:0] out1285; 
reg [127:0] out1286; 
reg [127:0] out1287; 
reg [127:0] out1288; 
reg [127:0] out1289; 
reg [127:0] out1290; 
reg [127:0] out1291; 
reg [127:0] out1292; 
reg [127:0] out1293; 
reg [127:0] out1294; 
reg [127:0] out1295; 
reg [127:0] out1296; 
reg [127:0] out1297; 
reg [127:0] out1298; 
reg [127:0] out1299; 
reg [127:0] out1300; 
reg [127:0] out1301; 
reg [127:0] out1302; 
reg [127:0] out1303; 
reg [127:0] out1304; 
reg [127:0] out1305; 
reg [127:0] out1306; 
reg [127:0] out1307; 
reg [127:0] out1308; 
reg [127:0] out1309; 
reg [127:0] out1310; 
reg [127:0] out1311; 
reg [127:0] out1312; 
reg [127:0] out1313; 
reg [127:0] out1314; 
reg [127:0] out1315; 
reg [127:0] out1316; 
reg [127:0] out1317; 
reg [127:0] out1318; 
reg [127:0] out1319; 
reg [127:0] out1320; 
reg [127:0] out1321; 
reg [127:0] out1322; 
reg [127:0] out1323; 
reg [127:0] out1324; 
reg [127:0] out1325; 
reg [127:0] out1326; 
reg [127:0] out1327; 
reg [127:0] out1328; 
reg [127:0] out1329; 
reg [127:0] out1330; 
reg [127:0] out1331; 
reg [127:0] out1332; 
reg [127:0] out1333; 
reg [127:0] out1334; 
reg [127:0] out1335; 
reg [127:0] out1336; 
reg [127:0] out1337; 
reg [127:0] out1338; 
reg [127:0] out1339; 
reg [127:0] out1340; 
reg [127:0] out1341; 
reg [127:0] out1342; 
reg [127:0] out1343; 
reg [127:0] out1344; 
reg [127:0] out1345; 
reg [127:0] out1346; 
reg [127:0] out1347; 
reg [127:0] out1348; 
reg [127:0] out1349; 
reg [127:0] out1350; 
reg [127:0] out1351; 
reg [127:0] out1352; 
reg [127:0] out1353; 
reg [127:0] out1354; 
reg [127:0] out1355; 
reg [127:0] out1356; 
reg [127:0] out1357; 
reg [127:0] out1358; 
reg [127:0] out1359; 
reg [127:0] out1360; 
reg [127:0] out1361; 
reg [127:0] out1362; 
reg [127:0] out1363; 
reg [127:0] out1364; 
reg [127:0] out1365; 
reg [127:0] out1366; 
reg [127:0] out1367; 
reg [127:0] out1368; 
reg [127:0] out1369; 
reg [127:0] out1370; 
reg [127:0] out1371; 
reg [127:0] out1372; 
reg [127:0] out1373; 
reg [127:0] out1374; 
reg [127:0] out1375; 
reg [127:0] out1376; 
reg [127:0] out1377; 
reg [127:0] out1378; 
reg [127:0] out1379; 
reg [127:0] out1380; 
reg [127:0] out1381; 
reg [127:0] out1382; 
reg [127:0] out1383; 
reg [127:0] out1384; 
reg [127:0] out1385; 
reg [127:0] out1386; 
reg [127:0] out1387; 
reg [127:0] out1388; 
reg [127:0] out1389; 
reg [127:0] out1390; 
reg [127:0] out1391; 
reg [127:0] out1392; 
reg [127:0] out1393; 
reg [127:0] out1394; 
reg [127:0] out1395; 
reg [127:0] out1396; 
reg [127:0] out1397; 
reg [127:0] out1398; 
reg [127:0] out1399; 
reg [127:0] out1400; 
reg [127:0] out1401; 
reg [127:0] out1402; 
reg [127:0] out1403; 
reg [127:0] out1404; 
reg [127:0] out1405; 
reg [127:0] out1406; 
reg [127:0] out1407; 
reg [127:0] out1408; 
reg [127:0] out1409; 
reg [127:0] out1410; 
reg [127:0] out1411; 
reg [127:0] out1412; 
reg [127:0] out1413; 
reg [127:0] out1414; 
reg [127:0] out1415; 
reg [127:0] out1416; 
reg [127:0] out1417; 
reg [127:0] out1418; 
reg [127:0] out1419; 
reg [127:0] out1420; 
reg [127:0] out1421; 
reg [127:0] out1422; 
reg [127:0] out1423; 
reg [127:0] out1424; 
reg [127:0] out1425; 
reg [127:0] out1426; 
reg [127:0] out1427; 
reg [127:0] out1428; 
reg [127:0] out1429; 
reg [127:0] out1430; 
reg [127:0] out1431; 
reg [127:0] out1432; 
reg [127:0] out1433; 
reg [127:0] out1434; 
reg [127:0] out1435; 
reg [127:0] out1436; 
reg [127:0] out1437; 
reg [127:0] out1438; 
reg [127:0] out1439; 
reg [127:0] out1440; 
reg [127:0] out1441; 
reg [127:0] out1442; 
reg [127:0] out1443; 
reg [127:0] out1444; 
reg [127:0] out1445; 
reg [127:0] out1446; 
reg [127:0] out1447; 
reg [127:0] out1448; 
reg [127:0] out1449; 
reg [127:0] out1450; 
reg [127:0] out1451; 
reg [127:0] out1452; 
reg [127:0] out1453; 
reg [127:0] out1454; 
reg [127:0] out1455; 
reg [127:0] out1456; 
reg [127:0] out1457; 
reg [127:0] out1458; 
reg [127:0] out1459; 
reg [127:0] out1460; 
reg [127:0] out1461; 
reg [127:0] out1462; 
reg [127:0] out1463; 
reg [127:0] out1464; 
reg [127:0] out1465; 
reg [127:0] out1466; 
reg [127:0] out1467; 
reg [127:0] out1468; 
reg [127:0] out1469; 
reg [127:0] out1470; 
reg [127:0] out1471; 
reg [127:0] out1472; 
reg [127:0] out1473; 
reg [127:0] out1474; 
reg [127:0] out1475; 
reg [127:0] out1476; 
reg [127:0] out1477; 
reg [127:0] out1478; 
reg [127:0] out1479; 
reg [127:0] out1480; 
reg [127:0] out1481; 
reg [127:0] out1482; 
reg [127:0] out1483; 
reg [127:0] out1484; 
reg [127:0] out1485; 
reg [127:0] out1486; 
reg [127:0] out1487; 
reg [127:0] out1488; 
reg [127:0] out1489; 
reg [127:0] out1490; 
reg [127:0] out1491; 
reg [127:0] out1492; 
reg [127:0] out1493; 
reg [127:0] out1494; 
reg [127:0] out1495; 
reg [127:0] out1496; 
reg [127:0] out1497; 
reg [127:0] out1498; 
reg [127:0] out1499; 
reg [127:0] out1500; 
reg [127:0] out1501; 
reg [127:0] out1502; 
reg [127:0] out1503; 
reg [127:0] out1504; 
reg [127:0] out1505; 
reg [127:0] out1506; 
reg [127:0] out1507; 
reg [127:0] out1508; 
reg [127:0] out1509; 
reg [127:0] out1510; 
reg [127:0] out1511; 
reg [127:0] out1512; 
reg [127:0] out1513; 
reg [127:0] out1514; 
reg [127:0] out1515; 
reg [127:0] out1516; 
reg [127:0] out1517; 
reg [127:0] out1518; 
reg [127:0] out1519; 
reg [127:0] out1520; 
reg [127:0] out1521; 
reg [127:0] out1522; 
reg [127:0] out1523; 
reg [127:0] out1524; 
reg [127:0] out1525; 
reg [127:0] out1526; 
reg [127:0] out1527; 
reg [127:0] out1528; 
reg [127:0] out1529; 
reg [127:0] out1530; 
reg [127:0] out1531; 
reg [127:0] out1532; 
reg [127:0] out1533; 
reg [127:0] out1534; 
reg [127:0] out1535; 
reg [127:0] out1536; 
reg [127:0] out1537; 
reg [127:0] out1538; 
reg [127:0] out1539; 
reg [127:0] out1540; 
reg [127:0] out1541; 
reg [127:0] out1542; 
reg [127:0] out1543; 
reg [127:0] out1544; 
reg [127:0] out1545; 
reg [127:0] out1546; 
reg [127:0] out1547; 
reg [127:0] out1548; 
reg [127:0] out1549; 
reg [127:0] out1550; 
reg [127:0] out1551; 
reg [127:0] out1552; 
reg [127:0] out1553; 
reg [127:0] out1554; 
reg [127:0] out1555; 
reg [127:0] out1556; 
reg [127:0] out1557; 
reg [127:0] out1558; 
reg [127:0] out1559; 
reg [127:0] out1560; 
reg [127:0] out1561; 
reg [127:0] out1562; 
reg [127:0] out1563; 
reg [127:0] out1564; 
reg [127:0] out1565; 
reg [127:0] out1566; 
reg [127:0] out1567; 
reg [127:0] out1568; 
reg [127:0] out1569; 
reg [127:0] out1570; 
reg [127:0] out1571; 
reg [127:0] out1572; 
reg [127:0] out1573; 
reg [127:0] out1574; 
reg [127:0] out1575; 
reg [127:0] out1576; 
reg [127:0] out1577; 
reg [127:0] out1578; 
reg [127:0] out1579; 
reg [127:0] out1580; 
reg [127:0] out1581; 
reg [127:0] out1582; 
reg [127:0] out1583; 
reg [127:0] out1584; 
reg [127:0] out1585; 
reg [127:0] out1586; 
reg [127:0] out1587; 
reg [127:0] out1588; 
reg [127:0] out1589; 
reg [127:0] out1590; 
reg [127:0] out1591; 
reg [127:0] out1592; 
reg [127:0] out1593; 
reg [127:0] out1594; 
reg [127:0] out1595; 
reg [127:0] out1596; 
reg [127:0] out1597; 
reg [127:0] out1598; 
reg [127:0] out1599; 
reg [127:0] out1600; 
reg [127:0] out1601; 
reg [127:0] out1602; 
reg [127:0] out1603; 
reg [127:0] out1604; 
reg [127:0] out1605; 
reg [127:0] out1606; 
reg [127:0] out1607; 
reg [127:0] out1608; 
reg [127:0] out1609; 
reg [127:0] out1610; 
reg [127:0] out1611; 
reg [127:0] out1612; 
reg [127:0] out1613; 
reg [127:0] out1614; 
reg [127:0] out1615; 
reg [127:0] out1616; 
reg [127:0] out1617; 
reg [127:0] out1618; 
reg [127:0] out1619; 
reg [127:0] out1620; 
reg [127:0] out1621; 
reg [127:0] out1622; 
reg [127:0] out1623; 
reg [127:0] out1624; 
reg [127:0] out1625; 
reg [127:0] out1626; 
reg [127:0] out1627; 
reg [127:0] out1628; 
reg [127:0] out1629; 
reg [127:0] out1630; 
reg [127:0] out1631; 
reg [127:0] out1632; 
reg [127:0] out1633; 
reg [127:0] out1634; 
reg [127:0] out1635; 
reg [127:0] out1636; 
reg [127:0] out1637; 
reg [127:0] out1638; 
reg [127:0] out1639; 
reg [127:0] out1640; 
reg [127:0] out1641; 
reg [127:0] out1642; 
reg [127:0] out1643; 
reg [127:0] out1644; 
reg [127:0] out1645; 
reg [127:0] out1646; 
reg [127:0] out1647; 
reg [127:0] out1648; 
reg [127:0] out1649; 
reg [127:0] out1650; 
reg [127:0] out1651; 
reg [127:0] out1652; 
reg [127:0] out1653; 
reg [127:0] out1654; 
reg [127:0] out1655; 
reg [127:0] out1656; 
reg [127:0] out1657; 
reg [127:0] out1658; 
reg [127:0] out1659; 
reg [127:0] out1660; 
reg [127:0] out1661; 
reg [127:0] out1662; 
reg [127:0] out1663; 
reg [127:0] out1664; 
reg [127:0] out1665; 
reg [127:0] out1666; 
reg [127:0] out1667; 
reg [127:0] out1668; 
reg [127:0] out1669; 
reg [127:0] out1670; 
reg [127:0] out1671; 
reg [127:0] out1672; 
reg [127:0] out1673; 
reg [127:0] out1674; 
reg [127:0] out1675; 
reg [127:0] out1676; 
reg [127:0] out1677; 
reg [127:0] out1678; 
reg [127:0] out1679; 
reg [127:0] out1680; 
reg [127:0] out1681; 
reg [127:0] out1682; 
reg [127:0] out1683; 
reg [127:0] out1684; 
reg [127:0] out1685; 
reg [127:0] out1686; 
reg [127:0] out1687; 
reg [127:0] out1688; 
reg [127:0] out1689; 
reg [127:0] out1690; 
reg [127:0] out1691; 
reg [127:0] out1692; 
reg [127:0] out1693; 
reg [127:0] out1694; 
reg [127:0] out1695; 
reg [127:0] out1696; 
reg [127:0] out1697; 
reg [127:0] out1698; 
reg [127:0] out1699; 
reg [127:0] out1700; 
reg [127:0] out1701; 
reg [127:0] out1702; 
reg [127:0] out1703; 
reg [127:0] out1704; 
reg [127:0] out1705; 
reg [127:0] out1706; 
reg [127:0] out1707; 
reg [127:0] out1708; 
reg [127:0] out1709; 
reg [127:0] out1710; 
reg [127:0] out1711; 
reg [127:0] out1712; 
reg [127:0] out1713; 
reg [127:0] out1714; 
reg [127:0] out1715; 
reg [127:0] out1716; 
reg [127:0] out1717; 
reg [127:0] out1718; 
reg [127:0] out1719; 
reg [127:0] out1720; 
reg [127:0] out1721; 
reg [127:0] out1722; 
reg [127:0] out1723; 
reg [127:0] out1724; 
reg [127:0] out1725; 
reg [127:0] out1726; 
reg [127:0] out1727; 
reg [127:0] out1728; 
reg [127:0] out1729; 
reg [127:0] out1730; 
reg [127:0] out1731; 
reg [127:0] out1732; 
reg [127:0] out1733; 
reg [127:0] out1734; 
reg [127:0] out1735; 
reg [127:0] out1736; 
reg [127:0] out1737; 
reg [127:0] out1738; 
reg [127:0] out1739; 
reg [127:0] out1740; 
reg [127:0] out1741; 
reg [127:0] out1742; 
reg [127:0] out1743; 
reg [127:0] out1744; 
reg [127:0] out1745; 
reg [127:0] out1746; 
reg [127:0] out1747; 
reg [127:0] out1748; 
reg [127:0] out1749; 
reg [127:0] out1750; 
reg [127:0] out1751; 
reg [127:0] out1752; 
reg [127:0] out1753; 
reg [127:0] out1754; 
reg [127:0] out1755; 
reg [127:0] out1756; 
reg [127:0] out1757; 
reg [127:0] out1758; 
reg [127:0] out1759; 
reg [127:0] out1760; 
reg [127:0] out1761; 
reg [127:0] out1762; 
reg [127:0] out1763; 
reg [127:0] out1764; 
reg [127:0] out1765; 
reg [127:0] out1766; 
reg [127:0] out1767; 
reg [127:0] out1768; 
reg [127:0] out1769; 
reg [127:0] out1770; 
reg [127:0] out1771; 
reg [127:0] out1772; 
reg [127:0] out1773; 
reg [127:0] out1774; 
reg [127:0] out1775; 
reg [127:0] out1776; 
reg [127:0] out1777; 
reg [127:0] out1778; 
reg [127:0] out1779; 
reg [127:0] out1780; 
reg [127:0] out1781; 
reg [127:0] out1782; 
reg [127:0] out1783; 
reg [127:0] out1784; 
reg [127:0] out1785; 
reg [127:0] out1786; 
reg [127:0] out1787; 
reg [127:0] out1788; 
reg [127:0] out1789; 
reg [127:0] out1790; 
reg [127:0] out1791; 
reg [127:0] out1792; 
reg [127:0] out1793; 
reg [127:0] out1794; 
reg [127:0] out1795; 
reg [127:0] out1796; 
reg [127:0] out1797; 
reg [127:0] out1798; 
reg [127:0] out1799; 
reg [127:0] out1800; 
reg [127:0] out1801; 
reg [127:0] out1802; 
reg [127:0] out1803; 
reg [127:0] out1804; 
reg [127:0] out1805; 
reg [127:0] out1806; 
reg [127:0] out1807; 
reg [127:0] out1808; 
reg [127:0] out1809; 
reg [127:0] out1810; 
reg [127:0] out1811; 
reg [127:0] out1812; 
reg [127:0] out1813; 
reg [127:0] out1814; 
reg [127:0] out1815; 
reg [127:0] out1816; 
reg [127:0] out1817; 
reg [127:0] out1818; 
reg [127:0] out1819; 
reg [127:0] out1820; 
reg [127:0] out1821; 
reg [127:0] out1822; 
reg [127:0] out1823; 
reg [127:0] out1824; 
reg [127:0] out1825; 
reg [127:0] out1826; 
reg [127:0] out1827; 
reg [127:0] out1828; 
reg [127:0] out1829; 
reg [127:0] out1830; 
reg [127:0] out1831; 
reg [127:0] out1832; 
reg [127:0] out1833; 
reg [127:0] out1834; 
reg [127:0] out1835; 
reg [127:0] out1836; 
reg [127:0] out1837; 
reg [127:0] out1838; 
reg [127:0] out1839; 
reg [127:0] out1840; 
reg [127:0] out1841; 
reg [127:0] out1842; 
reg [127:0] out1843; 
reg [127:0] out1844; 
reg [127:0] out1845; 
reg [127:0] out1846; 
reg [127:0] out1847; 
reg [127:0] out1848; 
reg [127:0] out1849; 
reg [127:0] out1850; 
reg [127:0] out1851; 
reg [127:0] out1852; 
reg [127:0] out1853; 
reg [127:0] out1854; 
reg [127:0] out1855; 
reg [127:0] out1856; 
reg [127:0] out1857; 
reg [127:0] out1858; 
reg [127:0] out1859; 
reg [127:0] out1860; 
reg [127:0] out1861; 
reg [127:0] out1862; 
reg [127:0] out1863; 
reg [127:0] out1864; 
reg [127:0] out1865; 
reg [127:0] out1866; 
reg [127:0] out1867; 
reg [127:0] out1868; 
reg [127:0] out1869; 
reg [127:0] out1870; 
reg [127:0] out1871; 
reg [127:0] out1872; 
reg [127:0] out1873; 
reg [127:0] out1874; 
reg [127:0] out1875; 
reg [127:0] out1876; 
reg [127:0] out1877; 
reg [127:0] out1878; 
reg [127:0] out1879; 
reg [127:0] out1880; 
reg [127:0] out1881; 
reg [127:0] out1882; 
reg [127:0] out1883; 
reg [127:0] out1884; 
reg [127:0] out1885; 
reg [127:0] out1886; 
reg [127:0] out1887; 
reg [127:0] out1888; 
reg [127:0] out1889; 
reg [127:0] out1890; 
reg [127:0] out1891; 
reg [127:0] out1892; 
reg [127:0] out1893; 
reg [127:0] out1894; 
reg [127:0] out1895; 
reg [127:0] out1896; 
reg [127:0] out1897; 
reg [127:0] out1898; 
reg [127:0] out1899; 
reg [127:0] out1900; 
reg [127:0] out1901; 
reg [127:0] out1902; 
reg [127:0] out1903; 
reg [127:0] out1904; 
reg [127:0] out1905; 
reg [127:0] out1906; 
reg [127:0] out1907; 
reg [127:0] out1908; 
reg [127:0] out1909; 
reg [127:0] out1910; 
reg [127:0] out1911; 
reg [127:0] out1912; 
reg [127:0] out1913; 
reg [127:0] out1914; 
reg [127:0] out1915; 
reg [127:0] out1916; 
reg [127:0] out1917; 
reg [127:0] out1918; 
reg [127:0] out1919; 
reg [127:0] out1920; 
reg [127:0] out1921; 
reg [127:0] out1922; 
reg [127:0] out1923; 
reg [127:0] out1924; 
reg [127:0] out1925; 
reg [127:0] out1926; 
reg [127:0] out1927; 
reg [127:0] out1928; 
reg [127:0] out1929; 
reg [127:0] out1930; 
reg [127:0] out1931; 
reg [127:0] out1932; 
reg [127:0] out1933; 
reg [127:0] out1934; 
reg [127:0] out1935; 
reg [127:0] out1936; 
reg [127:0] out1937; 
reg [127:0] out1938; 
reg [127:0] out1939; 
reg [127:0] out1940; 
reg [127:0] out1941; 
reg [127:0] out1942; 
reg [127:0] out1943; 
reg [127:0] out1944; 
reg [127:0] out1945; 
reg [127:0] out1946; 
reg [127:0] out1947; 
reg [127:0] out1948; 
reg [127:0] out1949; 
reg [127:0] out1950; 
reg [127:0] out1951; 
reg [127:0] out1952; 
reg [127:0] out1953; 
reg [127:0] out1954; 
reg [127:0] out1955; 
reg [127:0] out1956; 
reg [127:0] out1957; 
reg [127:0] out1958; 
reg [127:0] out1959; 
reg [127:0] out1960; 
reg [127:0] out1961; 
reg [127:0] out1962; 
reg [127:0] out1963; 
reg [127:0] out1964; 
reg [127:0] out1965; 
reg [127:0] out1966; 
reg [127:0] out1967; 
reg [127:0] out1968; 
reg [127:0] out1969; 
reg [127:0] out1970; 
reg [127:0] out1971; 
reg [127:0] out1972; 
reg [127:0] out1973; 
reg [127:0] out1974; 
reg [127:0] out1975; 
reg [127:0] out1976; 
reg [127:0] out1977; 
reg [127:0] out1978; 
reg [127:0] out1979; 
reg [127:0] out1980; 
reg [127:0] out1981; 
reg [127:0] out1982; 
reg [127:0] out1983; 
reg [127:0] out1984; 
reg [127:0] out1985; 
reg [127:0] out1986; 
reg [127:0] out1987; 
reg [127:0] out1988; 
reg [127:0] out1989; 
reg [127:0] out1990; 
reg [127:0] out1991; 
reg [127:0] out1992; 
reg [127:0] out1993; 
reg [127:0] out1994; 
reg [127:0] out1995; 
reg [127:0] out1996; 
reg [127:0] out1997; 
reg [127:0] out1998; 
reg [127:0] out1999; 
reg [127:0] out2000; 
reg [127:0] out2001; 
reg [127:0] out2002; 
reg [127:0] out2003; 
reg [127:0] out2004; 
reg [127:0] out2005; 
reg [127:0] out2006; 
reg [127:0] out2007; 
reg [127:0] out2008; 
reg [127:0] out2009; 
reg [127:0] out2010; 
reg [127:0] out2011; 
reg [127:0] out2012; 
reg [127:0] out2013; 
reg [127:0] out2014; 
reg [127:0] out2015; 
reg [127:0] out2016; 
reg [127:0] out2017; 
reg [127:0] out2018; 
reg [127:0] out2019; 
reg [127:0] out2020; 
reg [127:0] out2021; 
reg [127:0] out2022; 
reg [127:0] out2023; 
reg [127:0] out2024; 
reg [127:0] out2025; 
reg [127:0] out2026; 
reg [127:0] out2027; 
reg [127:0] out2028; 
reg [127:0] out2029; 
reg [127:0] out2030; 
reg [127:0] out2031; 
reg [127:0] out2032; 
reg [127:0] out2033; 
reg [127:0] out2034; 
reg [127:0] out2035; 
reg [127:0] out2036; 
reg [127:0] out2037; 
reg [127:0] out2038; 
reg [127:0] out2039; 
reg [127:0] out2040; 
reg [127:0] out2041; 
reg [127:0] out2042; 
reg [127:0] out2043; 
reg [127:0] out2044; 
reg [127:0] out2045; 
reg [127:0] out2046; 
reg [127:0] out2047; 
reg [127:0] out2048; 
reg [127:0] out2049; 
reg [127:0] out2050; 
reg [127:0] out2051; 
reg [127:0] out2052; 
reg [127:0] out2053; 
reg [127:0] out2054; 
reg [127:0] out2055; 
reg [127:0] out2056; 
reg [127:0] out2057; 
reg [127:0] out2058; 
reg [127:0] out2059; 
reg [127:0] out2060; 
reg [127:0] out2061; 
reg [127:0] out2062; 
reg [127:0] out2063; 
reg [127:0] out2064; 
reg [127:0] out2065; 
reg [127:0] out2066; 
reg [127:0] out2067; 
reg [127:0] out2068; 
reg [127:0] out2069; 
reg [127:0] out2070; 
reg [127:0] out2071; 
reg [127:0] out2072; 
reg [127:0] out2073; 
reg [127:0] out2074; 
reg [127:0] out2075; 
reg [127:0] out2076; 
reg [127:0] out2077; 
reg [127:0] out2078; 
reg [127:0] out2079; 
reg [127:0] out2080; 
reg [127:0] out2081; 
reg [127:0] out2082; 
reg [127:0] out2083; 
reg [127:0] out2084; 
reg [127:0] out2085; 
reg [127:0] out2086; 
reg [127:0] out2087; 
reg [127:0] out2088; 
reg [127:0] out2089; 
reg [127:0] out2090; 
reg [127:0] out2091; 
reg [127:0] out2092; 
reg [127:0] out2093; 
reg [127:0] out2094; 
reg [127:0] out2095; 
reg [127:0] out2096; 
reg [127:0] out2097; 
reg [127:0] out2098; 
reg [127:0] out2099; 
reg [127:0] out2100; 
reg [127:0] out2101; 
reg [127:0] out2102; 
reg [127:0] out2103; 
reg [127:0] out2104; 
reg [127:0] out2105; 
reg [127:0] out2106; 
reg [127:0] out2107; 
reg [127:0] out2108; 
reg [127:0] out2109; 
reg [127:0] out2110; 
reg [127:0] out2111; 
reg [127:0] out2112; 
reg [127:0] out2113; 
reg [127:0] out2114; 
reg [127:0] out2115; 
reg [127:0] out2116; 
reg [127:0] out2117; 
reg [127:0] out2118; 
reg [127:0] out2119; 
reg [127:0] out2120; 
reg [127:0] out2121; 
reg [127:0] out2122; 
reg [127:0] out2123; 
reg [127:0] out2124; 
reg [127:0] out2125; 
reg [127:0] out2126; 
reg [127:0] out2127; 
reg [127:0] out2128; 
reg [127:0] out2129; 
reg [127:0] out2130; 
reg [127:0] out2131; 
reg [127:0] out2132; 
reg [127:0] out2133; 
reg [127:0] out2134; 
reg [127:0] out2135; 
reg [127:0] out2136; 
reg [127:0] out2137; 
reg [127:0] out2138; 
reg [127:0] out2139; 
reg [127:0] out2140; 
reg [127:0] out2141; 
reg [127:0] out2142; 
reg [127:0] out2143; 
reg [127:0] out2144; 
reg [127:0] out2145; 
reg [127:0] out2146; 
reg [127:0] out2147; 
reg [127:0] out2148; 
reg [127:0] out2149; 
reg [127:0] out2150; 
reg [127:0] out2151; 
reg [127:0] out2152; 
reg [127:0] out2153; 
reg [127:0] out2154; 
reg [127:0] out2155; 
reg [127:0] out2156; 
reg [127:0] out2157; 
reg [127:0] out2158; 
reg [127:0] out2159; 
reg [127:0] out2160; 
reg [127:0] out2161; 
reg [127:0] out2162; 
reg [127:0] out2163; 
reg [127:0] out2164; 
reg [127:0] out2165; 
reg [127:0] out2166; 
reg [127:0] out2167; 
reg [127:0] out2168; 
reg [127:0] out2169; 
reg [127:0] out2170; 
reg [127:0] out2171; 
reg [127:0] out2172; 
reg [127:0] out2173; 
reg [127:0] out2174; 
reg [127:0] out2175; 
reg [127:0] out2176; 
reg [127:0] out2177; 
reg [127:0] out2178; 
reg [127:0] out2179; 
reg [127:0] out2180; 
reg [127:0] out2181; 
reg [127:0] out2182; 
reg [127:0] out2183; 
reg [127:0] out2184; 
reg [127:0] out2185; 
reg [127:0] out2186; 
reg [127:0] out2187; 
reg [127:0] out2188; 
reg [127:0] out2189; 
reg [127:0] out2190; 
reg [127:0] out2191; 
reg [127:0] out2192; 
reg [127:0] out2193; 
reg [127:0] out2194; 
reg [127:0] out2195; 
reg [127:0] out2196; 
reg [127:0] out2197; 
reg [127:0] out2198; 
reg [127:0] out2199; 
reg [127:0] out2200; 
reg [127:0] out2201; 
reg [127:0] out2202; 
reg [127:0] out2203; 
reg [127:0] out2204; 
reg [127:0] out2205; 
reg [127:0] out2206; 
reg [127:0] out2207; 
reg [127:0] out2208; 
reg [127:0] out2209; 
reg [127:0] out2210; 
reg [127:0] out2211; 
reg [127:0] out2212; 
reg [127:0] out2213; 
reg [127:0] out2214; 
reg [127:0] out2215; 
reg [127:0] out2216; 
reg [127:0] out2217; 
reg [127:0] out2218; 
reg [127:0] out2219; 
reg [127:0] out2220; 
reg [127:0] out2221; 
reg [127:0] out2222; 
reg [127:0] out2223; 
reg [127:0] out2224; 
reg [127:0] out2225; 
reg [127:0] out2226; 
reg [127:0] out2227; 
reg [127:0] out2228; 
reg [127:0] out2229; 
reg [127:0] out2230; 
reg [127:0] out2231; 
reg [127:0] out2232; 
reg [127:0] out2233; 
reg [127:0] out2234; 
reg [127:0] out2235; 
reg [127:0] out2236; 
reg [127:0] out2237; 
reg [127:0] out2238; 
reg [127:0] out2239; 
reg [127:0] out2240; 
reg [127:0] out2241; 
reg [127:0] out2242; 
reg [127:0] out2243; 
reg [127:0] out2244; 
reg [127:0] out2245; 
reg [127:0] out2246; 
reg [127:0] out2247; 
reg [127:0] out2248; 
reg [127:0] out2249; 
reg [127:0] out2250; 
reg [127:0] out2251; 
reg [127:0] out2252; 
reg [127:0] out2253; 
reg [127:0] out2254; 
reg [127:0] out2255; 
reg [127:0] out2256; 
reg [127:0] out2257; 
reg [127:0] out2258; 
reg [127:0] out2259; 
reg [127:0] out2260; 
reg [127:0] out2261; 
reg [127:0] out2262; 
reg [127:0] out2263; 
reg [127:0] out2264; 
reg [127:0] out2265; 
reg [127:0] out2266; 
reg [127:0] out2267; 
reg [127:0] out2268; 
reg [127:0] out2269; 
reg [127:0] out2270; 
reg [127:0] out2271; 
reg [127:0] out2272; 
reg [127:0] out2273; 
reg [127:0] out2274; 
reg [127:0] out2275; 
reg [127:0] out2276; 
reg [127:0] out2277; 
reg [127:0] out2278; 
reg [127:0] out2279; 
reg [127:0] out2280; 
reg [127:0] out2281; 
reg [127:0] out2282; 
reg [127:0] out2283; 
reg [127:0] out2284; 
reg [127:0] out2285; 
reg [127:0] out2286; 
reg [127:0] out2287; 
reg [127:0] out2288; 
reg [127:0] out2289; 
reg [127:0] out2290; 
reg [127:0] out2291; 
reg [127:0] out2292; 
reg [127:0] out2293; 
reg [127:0] out2294; 
reg [127:0] out2295; 
reg [127:0] out2296; 
reg [127:0] out2297; 
reg [127:0] out2298; 
reg [127:0] out2299; 
reg [127:0] out2300; 
reg [127:0] out2301; 
reg [127:0] out2302; 
reg [127:0] out2303; 
reg [127:0] out2304; 
reg [127:0] out2305; 
reg [127:0] out2306; 
reg [127:0] out2307; 
reg [127:0] out2308; 
reg [127:0] out2309; 
reg [127:0] out2310; 
reg [127:0] out2311; 
reg [127:0] out2312; 
reg [127:0] out2313; 
reg [127:0] out2314; 
reg [127:0] out2315; 
reg [127:0] out2316; 
reg [127:0] out2317; 
reg [127:0] out2318; 
reg [127:0] out2319; 
reg [127:0] out2320; 
reg [127:0] out2321; 
reg [127:0] out2322; 
reg [127:0] out2323; 
reg [127:0] out2324; 
reg [127:0] out2325; 
reg [127:0] out2326; 
reg [127:0] out2327; 
reg [127:0] out2328; 
reg [127:0] out2329; 
reg [127:0] out2330; 
reg [127:0] out2331; 
reg [127:0] out2332; 
reg [127:0] out2333; 
reg [127:0] out2334; 
reg [127:0] out2335; 
reg [127:0] out2336; 
reg [127:0] out2337; 
reg [127:0] out2338; 
reg [127:0] out2339; 
reg [127:0] out2340; 
reg [127:0] out2341; 
reg [127:0] out2342; 
reg [127:0] out2343; 
reg [127:0] out2344; 
reg [127:0] out2345; 
reg [127:0] out2346; 
reg [127:0] out2347; 
reg [127:0] out2348; 
reg [127:0] out2349; 
reg [127:0] out2350; 
reg [127:0] out2351; 
reg [127:0] out2352; 
reg [127:0] out2353; 
reg [127:0] out2354; 
reg [127:0] out2355; 
reg [127:0] out2356; 
reg [127:0] out2357; 
reg [127:0] out2358; 
reg [127:0] out2359; 
reg [127:0] out2360; 
reg [127:0] out2361; 
reg [127:0] out2362; 
reg [127:0] out2363; 
reg [127:0] out2364; 
reg [127:0] out2365; 
reg [127:0] out2366; 
reg [127:0] out2367; 
reg [127:0] out2368; 
reg [127:0] out2369; 
reg [127:0] out2370; 
reg [127:0] out2371; 
reg [127:0] out2372; 
reg [127:0] out2373; 
reg [127:0] out2374; 
reg [127:0] out2375; 
reg [127:0] out2376; 
reg [127:0] out2377; 
reg [127:0] out2378; 
reg [127:0] out2379; 
reg [127:0] out2380; 
reg [127:0] out2381; 
reg [127:0] out2382; 
reg [127:0] out2383; 
reg [127:0] out2384; 
reg [127:0] out2385; 
reg [127:0] out2386; 
reg [127:0] out2387; 
reg [127:0] out2388; 
reg [127:0] out2389; 
reg [127:0] out2390; 
reg [127:0] out2391; 
reg [127:0] out2392; 
reg [127:0] out2393; 
reg [127:0] out2394; 
reg [127:0] out2395; 
reg [127:0] out2396; 
reg [127:0] out2397; 
reg [127:0] out2398; 
reg [127:0] out2399; 
reg [127:0] out2400; 
reg [127:0] out2401; 
reg [127:0] out2402; 
reg [127:0] out2403; 
reg [127:0] out2404; 
reg [127:0] out2405; 
reg [127:0] out2406; 
reg [127:0] out2407; 
reg [127:0] out2408; 
reg [127:0] out2409; 
reg [127:0] out2410; 
reg [127:0] out2411; 
reg [127:0] out2412; 
reg [127:0] out2413; 
reg [127:0] out2414; 
reg [127:0] out2415; 
reg [127:0] out2416; 
reg [127:0] out2417; 
reg [127:0] out2418; 
reg [127:0] out2419; 
reg [127:0] out2420; 
reg [127:0] out2421; 
reg [127:0] out2422; 
reg [127:0] out2423; 
reg [127:0] out2424; 
reg [127:0] out2425; 
reg [127:0] out2426; 
reg [127:0] out2427; 
reg [127:0] out2428; 
reg [127:0] out2429; 
reg [127:0] out2430; 
reg [127:0] out2431; 
reg [127:0] out2432; 
reg [127:0] out2433; 
reg [127:0] out2434; 
reg [127:0] out2435; 
reg [127:0] out2436; 
reg [127:0] out2437; 
reg [127:0] out2438; 
reg [127:0] out2439; 
reg [127:0] out2440; 
reg [127:0] out2441; 
reg [127:0] out2442; 
reg [127:0] out2443; 
reg [127:0] out2444; 
reg [127:0] out2445; 
reg [127:0] out2446; 
reg [127:0] out2447; 
reg [127:0] out2448; 
reg [127:0] out2449; 
reg [127:0] out2450; 
reg [127:0] out2451; 
reg [127:0] out2452; 
reg [127:0] out2453; 
reg [127:0] out2454; 
reg [127:0] out2455; 
reg [127:0] out2456; 
reg [127:0] out2457; 
reg [127:0] out2458; 
reg [127:0] out2459; 
reg [127:0] out2460; 
reg [127:0] out2461; 
reg [127:0] out2462; 
reg [127:0] out2463; 
reg [127:0] out2464; 
reg [127:0] out2465; 
reg [127:0] out2466; 
reg [127:0] out2467; 
reg [127:0] out2468; 
reg [127:0] out2469; 
reg [127:0] out2470; 
reg [127:0] out2471; 
reg [127:0] out2472; 
reg [127:0] out2473; 
reg [127:0] out2474; 
reg [127:0] out2475; 
reg [127:0] out2476; 
reg [127:0] out2477; 
reg [127:0] out2478; 
reg [127:0] out2479; 
reg [127:0] out2480; 
reg [127:0] out2481; 
reg [127:0] out2482; 
reg [127:0] out2483; 
reg [127:0] out2484; 
reg [127:0] out2485; 
reg [127:0] out2486; 
reg [127:0] out2487; 
reg [127:0] out2488; 
reg [127:0] out2489; 
reg [127:0] out2490; 
reg [127:0] out2491; 
reg [127:0] out2492; 
reg [127:0] out2493; 
reg [127:0] out2494; 
reg [127:0] out2495; 
reg [127:0] out2496; 
reg [127:0] out2497; 
reg [127:0] out2498; 
reg [127:0] out2499; 
reg [127:0] out2500; 
reg [127:0] out2501; 
reg [127:0] out2502; 
reg [127:0] out2503; 
reg [127:0] out2504; 
reg [127:0] out2505; 
reg [127:0] out2506; 
reg [127:0] out2507; 
reg [127:0] out2508; 
reg [127:0] out2509; 
reg [127:0] out2510; 
reg [127:0] out2511; 
reg [127:0] out2512; 
reg [127:0] out2513; 
reg [127:0] out2514; 
reg [127:0] out2515; 
reg [127:0] out2516; 
reg [127:0] out2517; 
reg [127:0] out2518; 
reg [127:0] out2519; 
reg [127:0] out2520; 
reg [127:0] out2521; 
reg [127:0] out2522; 
reg [127:0] out2523; 
reg [127:0] out2524; 
reg [127:0] out2525; 
reg [127:0] out2526; 
reg [127:0] out2527; 
reg [127:0] out2528; 
reg [127:0] out2529; 
reg [127:0] out2530; 
reg [127:0] out2531; 
reg [127:0] out2532; 
reg [127:0] out2533; 
reg [127:0] out2534; 
reg [127:0] out2535; 
reg [127:0] out2536; 
reg [127:0] out2537; 
reg [127:0] out2538; 
reg [127:0] out2539; 
reg [127:0] out2540; 
reg [127:0] out2541; 
reg [127:0] out2542; 
reg [127:0] out2543; 
reg [127:0] out2544; 
reg [127:0] out2545; 
reg [127:0] out2546; 
reg [127:0] out2547; 
reg [127:0] out2548; 
reg [127:0] out2549; 
reg [127:0] out2550; 
reg [127:0] out2551; 
reg [127:0] out2552; 
reg [127:0] out2553; 
reg [127:0] out2554; 
reg [127:0] out2555; 
reg [127:0] out2556; 
reg [127:0] out2557; 
reg [127:0] out2558; 
reg [127:0] out2559; 
reg [127:0] out2560; 
reg [127:0] out2561; 
reg [127:0] out2562; 
reg [127:0] out2563; 
reg [127:0] out2564; 
reg [127:0] out2565; 
reg [127:0] out2566; 
reg [127:0] out2567; 
reg [127:0] out2568; 
reg [127:0] out2569; 
reg [127:0] out2570; 
reg [127:0] out2571; 
reg [127:0] out2572; 
reg [127:0] out2573; 
reg [127:0] out2574; 
reg [127:0] out2575; 
reg [127:0] out2576; 
reg [127:0] out2577; 
reg [127:0] out2578; 
reg [127:0] out2579; 
reg [127:0] out2580; 
reg [127:0] out2581; 
reg [127:0] out2582; 
reg [127:0] out2583; 
reg [127:0] out2584; 
reg [127:0] out2585; 
reg [127:0] out2586; 
reg [127:0] out2587; 
reg [127:0] out2588; 
reg [127:0] out2589; 
reg [127:0] out2590; 
reg [127:0] out2591; 
reg [127:0] out2592; 
reg [127:0] out2593; 
reg [127:0] out2594; 
reg [127:0] out2595; 
reg [127:0] out2596; 
reg [127:0] out2597; 
reg [127:0] out2598; 
reg [127:0] out2599; 
reg [127:0] out2600; 
reg [127:0] out2601; 
reg [127:0] out2602; 
reg [127:0] out2603; 
reg [127:0] out2604; 
reg [127:0] out2605; 
reg [127:0] out2606; 
reg [127:0] out2607; 
reg [127:0] out2608; 
reg [127:0] out2609; 
reg [127:0] out2610; 
reg [127:0] out2611; 
reg [127:0] out2612; 
reg [127:0] out2613; 
reg [127:0] out2614; 
reg [127:0] out2615; 
reg [127:0] out2616; 
reg [127:0] out2617; 
reg [127:0] out2618; 
reg [127:0] out2619; 
reg [127:0] out2620; 
reg [127:0] out2621; 
reg [127:0] out2622; 
reg [127:0] out2623; 
reg [127:0] out2624; 
reg [127:0] out2625; 
reg [127:0] out2626; 
reg [127:0] out2627; 
reg [127:0] out2628; 
reg [127:0] out2629; 
reg [127:0] out2630; 
reg [127:0] out2631; 
reg [127:0] out2632; 
reg [127:0] out2633; 
reg [127:0] out2634; 
reg [127:0] out2635; 
reg [127:0] out2636; 
reg [127:0] out2637; 
reg [127:0] out2638; 
reg [127:0] out2639; 
reg [127:0] out2640; 
reg [127:0] out2641; 
reg [127:0] out2642; 
reg [127:0] out2643; 
reg [127:0] out2644; 
reg [127:0] out2645; 
reg [127:0] out2646; 
reg [127:0] out2647; 
reg [127:0] out2648; 
reg [127:0] out2649; 
reg [127:0] out2650; 
reg [127:0] out2651; 
reg [127:0] out2652; 
reg [127:0] out2653; 
reg [127:0] out2654; 
reg [127:0] out2655; 
reg [127:0] out2656; 
reg [127:0] out2657; 
reg [127:0] out2658; 
reg [127:0] out2659; 
reg [127:0] out2660; 
reg [127:0] out2661; 
reg [127:0] out2662; 
reg [127:0] out2663; 
reg [127:0] out2664; 
reg [127:0] out2665; 
reg [127:0] out2666; 
reg [127:0] out2667; 
reg [127:0] out2668; 
reg [127:0] out2669; 
reg [127:0] out2670; 
reg [127:0] out2671; 
reg [127:0] out2672; 
reg [127:0] out2673; 
reg [127:0] out2674; 
reg [127:0] out2675; 
reg [127:0] out2676; 
reg [127:0] out2677; 
reg [127:0] out2678; 
reg [127:0] out2679; 
reg [127:0] out2680; 
reg [127:0] out2681; 
reg [127:0] out2682; 
reg [127:0] out2683; 
reg [127:0] out2684; 
reg [127:0] out2685; 
reg [127:0] out2686; 
reg [127:0] out2687; 
reg [127:0] out2688; 
reg [127:0] out2689; 
reg [127:0] out2690; 
reg [127:0] out2691; 
reg [127:0] out2692; 
reg [127:0] out2693; 
reg [127:0] out2694; 
reg [127:0] out2695; 
reg [127:0] out2696; 
reg [127:0] out2697; 
reg [127:0] out2698; 
reg [127:0] out2699; 
reg [127:0] out2700; 
reg [127:0] out2701; 
reg [127:0] out2702; 
reg [127:0] out2703; 
reg [127:0] out2704; 
reg [127:0] out2705; 
reg [127:0] out2706; 
reg [127:0] out2707; 
reg [127:0] out2708; 
reg [127:0] out2709; 
reg [127:0] out2710; 
reg [127:0] out2711; 
reg [127:0] out2712; 
reg [127:0] out2713; 
reg [127:0] out2714; 
reg [127:0] out2715; 
reg [127:0] out2716; 
reg [127:0] out2717; 
reg [127:0] out2718; 
reg [127:0] out2719; 
reg [127:0] out2720; 
reg [127:0] out2721; 
reg [127:0] out2722; 
reg [127:0] out2723; 
reg [127:0] out2724; 
reg [127:0] out2725; 
reg [127:0] out2726; 
reg [127:0] out2727; 
reg [127:0] out2728; 
reg [127:0] out2729; 
reg [127:0] out2730; 
reg [127:0] out2731; 
reg [127:0] out2732; 
reg [127:0] out2733; 
reg [127:0] out2734; 
reg [127:0] out2735; 
reg [127:0] out2736; 
reg [127:0] out2737; 
reg [127:0] out2738; 
reg [127:0] out2739; 
reg [127:0] out2740; 
reg [127:0] out2741; 
reg [127:0] out2742; 
reg [127:0] out2743; 
reg [127:0] out2744; 
reg [127:0] out2745; 
reg [127:0] out2746; 
reg [127:0] out2747; 
reg [127:0] out2748; 
reg [127:0] out2749; 
reg [127:0] out2750; 
reg [127:0] out2751; 
reg [127:0] out2752; 
reg [127:0] out2753; 
reg [127:0] out2754; 
reg [127:0] out2755; 
reg [127:0] out2756; 
reg [127:0] out2757; 
reg [127:0] out2758; 
reg [127:0] out2759; 
reg [127:0] out2760; 
reg [127:0] out2761; 
reg [127:0] out2762; 
reg [127:0] out2763; 
reg [127:0] out2764; 
reg [127:0] out2765; 
reg [127:0] out2766; 
reg [127:0] out2767; 
reg [127:0] out2768; 
reg [127:0] out2769; 
reg [127:0] out2770; 
reg [127:0] out2771; 
reg [127:0] out2772; 
reg [127:0] out2773; 
reg [127:0] out2774; 
reg [127:0] out2775; 
reg [127:0] out2776; 
reg [127:0] out2777; 
reg [127:0] out2778; 
reg [127:0] out2779; 
reg [127:0] out2780; 
reg [127:0] out2781; 
reg [127:0] out2782; 
reg [127:0] out2783; 
reg [127:0] out2784; 
reg [127:0] out2785; 
reg [127:0] out2786; 
reg [127:0] out2787; 
reg [127:0] out2788; 
reg [127:0] out2789; 
reg [127:0] out2790; 
reg [127:0] out2791; 
reg [127:0] out2792; 
reg [127:0] out2793; 
reg [127:0] out2794; 
reg [127:0] out2795; 
reg [127:0] out2796; 
reg [127:0] out2797; 
reg [127:0] out2798; 
reg [127:0] out2799; 
reg [127:0] out2800; 
reg [127:0] out2801; 
reg [127:0] out2802; 
reg [127:0] out2803; 
reg [127:0] out2804; 
reg [127:0] out2805; 
reg [127:0] out2806; 
reg [127:0] out2807; 
reg [127:0] out2808; 
reg [127:0] out2809; 
reg [127:0] out2810; 
reg [127:0] out2811; 
reg [127:0] out2812; 
reg [127:0] out2813; 
reg [127:0] out2814; 
reg [127:0] out2815; 
reg [127:0] out2816; 
reg [127:0] out2817; 
reg [127:0] out2818; 
reg [127:0] out2819; 
reg [127:0] out2820; 
reg [127:0] out2821; 
reg [127:0] out2822; 
reg [127:0] out2823; 
reg [127:0] out2824; 
reg [127:0] out2825; 
reg [127:0] out2826; 
reg [127:0] out2827; 
reg [127:0] out2828; 
reg [127:0] out2829; 
reg [127:0] out2830; 
reg [127:0] out2831; 
reg [127:0] out2832; 
reg [127:0] out2833; 
reg [127:0] out2834; 
reg [127:0] out2835; 
reg [127:0] out2836; 
reg [127:0] out2837; 
reg [127:0] out2838; 
reg [127:0] out2839; 
reg [127:0] out2840; 
reg [127:0] out2841; 
reg [127:0] out2842; 
reg [127:0] out2843; 
reg [127:0] out2844; 
reg [127:0] out2845; 
reg [127:0] out2846; 
reg [127:0] out2847; 
reg [127:0] out2848; 
reg [127:0] out2849; 
reg [127:0] out2850; 
reg [127:0] out2851; 
reg [127:0] out2852; 
reg [127:0] out2853; 
reg [127:0] out2854; 
reg [127:0] out2855; 
reg [127:0] out2856; 
reg [127:0] out2857; 
reg [127:0] out2858; 
reg [127:0] out2859; 
reg [127:0] out2860; 
reg [127:0] out2861; 
reg [127:0] out2862; 
reg [127:0] out2863; 
reg [127:0] out2864; 
reg [127:0] out2865; 
reg [127:0] out2866; 
reg [127:0] out2867; 
reg [127:0] out2868; 
reg [127:0] out2869; 
reg [127:0] out2870; 
reg [127:0] out2871; 
reg [127:0] out2872; 
reg [127:0] out2873; 
reg [127:0] out2874; 
reg [127:0] out2875; 
reg [127:0] out2876; 
reg [127:0] out2877; 
reg [127:0] out2878; 
reg [127:0] out2879; 
reg [127:0] out2880; 
reg [127:0] out2881; 
reg [127:0] out2882; 
reg [127:0] out2883; 
reg [127:0] out2884; 
reg [127:0] out2885; 
reg [127:0] out2886; 
reg [127:0] out2887; 
reg [127:0] out2888; 
reg [127:0] out2889; 
reg [127:0] out2890; 
reg [127:0] out2891; 
reg [127:0] out2892; 
reg [127:0] out2893; 
reg [127:0] out2894; 
reg [127:0] out2895; 
reg [127:0] out2896; 
reg [127:0] out2897; 
reg [127:0] out2898; 
reg [127:0] out2899; 
reg [127:0] out2900; 
reg [127:0] out2901; 
reg [127:0] out2902; 
reg [127:0] out2903; 
reg [127:0] out2904; 
reg [127:0] out2905; 
reg [127:0] out2906; 
reg [127:0] out2907; 
reg [127:0] out2908; 
reg [127:0] out2909; 
reg [127:0] out2910; 
reg [127:0] out2911; 
reg [127:0] out2912; 
reg [127:0] out2913; 
reg [127:0] out2914; 
reg [127:0] out2915; 
reg [127:0] out2916; 
reg [127:0] out2917; 
reg [127:0] out2918; 
reg [127:0] out2919; 
reg [127:0] out2920; 
reg [127:0] out2921; 
reg [127:0] out2922; 
reg [127:0] out2923; 
reg [127:0] out2924; 
reg [127:0] out2925; 
reg [127:0] out2926; 
reg [127:0] out2927; 
reg [127:0] out2928; 
reg [127:0] out2929; 
reg [127:0] out2930; 
reg [127:0] out2931; 
reg [127:0] out2932; 
reg [127:0] out2933; 
reg [127:0] out2934; 
reg [127:0] out2935; 
reg [127:0] out2936; 
reg [127:0] out2937; 
reg [127:0] out2938; 
reg [127:0] out2939; 
reg [127:0] out2940; 
reg [127:0] out2941; 
reg [127:0] out2942; 
reg [127:0] out2943; 
reg [127:0] out2944; 
reg [127:0] out2945; 
reg [127:0] out2946; 
reg [127:0] out2947; 
reg [127:0] out2948; 
reg [127:0] out2949; 
reg [127:0] out2950; 
reg [127:0] out2951; 
reg [127:0] out2952; 
reg [127:0] out2953; 
reg [127:0] out2954; 
reg [127:0] out2955; 
reg [127:0] out2956; 
reg [127:0] out2957; 
reg [127:0] out2958; 
reg [127:0] out2959; 
reg [127:0] out2960; 
reg [127:0] out2961; 
reg [127:0] out2962; 
reg [127:0] out2963; 
reg [127:0] out2964; 
reg [127:0] out2965; 
reg [127:0] out2966; 
reg [127:0] out2967; 
reg [127:0] out2968; 
reg [127:0] out2969; 
reg [127:0] out2970; 
reg [127:0] out2971; 
reg [127:0] out2972; 
reg [127:0] out2973; 
reg [127:0] out2974; 
reg [127:0] out2975; 
reg [127:0] out2976; 
reg [127:0] out2977; 
reg [127:0] out2978; 
reg [127:0] out2979; 
reg [127:0] out2980; 
reg [127:0] out2981; 
reg [127:0] out2982; 
reg [127:0] out2983; 
reg [127:0] out2984; 
reg [127:0] out2985; 
reg [127:0] out2986; 
reg [127:0] out2987; 
reg [127:0] out2988; 
reg [127:0] out2989; 
reg [127:0] out2990; 
reg [127:0] out2991; 
reg [127:0] out2992; 
reg [127:0] out2993; 
reg [127:0] out2994; 
reg [127:0] out2995; 
reg [127:0] out2996; 
reg [127:0] out2997; 
reg [127:0] out2998; 
reg [127:0] out2999; 
reg [127:0] out3000; 
reg [127:0] out3001; 
reg [127:0] out3002; 
reg [127:0] out3003; 
reg [127:0] out3004; 
reg [127:0] out3005; 
reg [127:0] out3006; 
reg [127:0] out3007; 
reg [127:0] out3008; 
reg [127:0] out3009; 
reg [127:0] out3010; 
reg [127:0] out3011; 
reg [127:0] out3012; 
reg [127:0] out3013; 
reg [127:0] out3014; 
reg [127:0] out3015; 
reg [127:0] out3016; 
reg [127:0] out3017; 
reg [127:0] out3018; 
reg [127:0] out3019; 
reg [127:0] out3020; 
reg [127:0] out3021; 
reg [127:0] out3022; 
reg [127:0] out3023; 
reg [127:0] out3024; 
reg [127:0] out3025; 
reg [127:0] out3026; 
reg [127:0] out3027; 
reg [127:0] out3028; 
reg [127:0] out3029; 
reg [127:0] out3030; 
reg [127:0] out3031; 
reg [127:0] out3032; 
reg [127:0] out3033; 
reg [127:0] out3034; 
reg [127:0] out3035; 
reg [127:0] out3036; 
reg [127:0] out3037; 
reg [127:0] out3038; 
reg [127:0] out3039; 
reg [127:0] out3040; 
reg [127:0] out3041; 
reg [127:0] out3042; 
reg [127:0] out3043; 
reg [127:0] out3044; 
reg [127:0] out3045; 
reg [127:0] out3046; 
reg [127:0] out3047; 
reg [127:0] out3048; 
reg [127:0] out3049; 
reg [127:0] out3050; 
reg [127:0] out3051; 
reg [127:0] out3052; 
reg [127:0] out3053; 
reg [127:0] out3054; 
reg [127:0] out3055; 
reg [127:0] out3056; 
reg [127:0] out3057; 
reg [127:0] out3058; 
reg [127:0] out3059; 
reg [127:0] out3060; 
reg [127:0] out3061; 
reg [127:0] out3062; 
reg [127:0] out3063; 
reg [127:0] out3064; 
reg [127:0] out3065; 
reg [127:0] out3066; 
reg [127:0] out3067; 
reg [127:0] out3068; 
reg [127:0] out3069; 
reg [127:0] out3070; 
reg [127:0] out3071; 
reg [127:0] out3072; 
reg [127:0] out3073; 
reg [127:0] out3074; 
reg [127:0] out3075; 
reg [127:0] out3076; 
reg [127:0] out3077; 
reg [127:0] out3078; 
reg [127:0] out3079; 
reg [127:0] out3080; 
reg [127:0] out3081; 
reg [127:0] out3082; 
reg [127:0] out3083; 
reg [127:0] out3084; 
reg [127:0] out3085; 
reg [127:0] out3086; 
reg [127:0] out3087; 
reg [127:0] out3088; 
reg [127:0] out3089; 
reg [127:0] out3090; 
reg [127:0] out3091; 
reg [127:0] out3092; 
reg [127:0] out3093; 
reg [127:0] out3094; 
reg [127:0] out3095; 
reg [127:0] out3096; 
reg [127:0] out3097; 
reg [127:0] out3098; 
reg [127:0] out3099; 
reg [127:0] out3100; 
reg [127:0] out3101; 
reg [127:0] out3102; 
reg [127:0] out3103; 
reg [127:0] out3104; 
reg [127:0] out3105; 
reg [127:0] out3106; 
reg [127:0] out3107; 
reg [127:0] out3108; 
reg [127:0] out3109; 
reg [127:0] out3110; 
reg [127:0] out3111; 
reg [127:0] out3112; 
reg [127:0] out3113; 
reg [127:0] out3114; 
reg [127:0] out3115; 
reg [127:0] out3116; 
reg [127:0] out3117; 
reg [127:0] out3118; 
reg [127:0] out3119; 
reg [127:0] out3120; 
reg [127:0] out3121; 
reg [127:0] out3122; 
reg [127:0] out3123; 
reg [127:0] out3124; 
reg [127:0] out3125; 
reg [127:0] out3126; 
reg [127:0] out3127; 
reg [127:0] out3128; 
reg [127:0] out3129; 
reg [127:0] out3130; 
reg [127:0] out3131; 
reg [127:0] out3132; 
reg [127:0] out3133; 
reg [127:0] out3134; 
reg [127:0] out3135; 
reg [127:0] out3136; 
reg [127:0] out3137; 
reg [127:0] out3138; 
reg [127:0] out3139; 
reg [127:0] out3140; 
reg [127:0] out3141; 
reg [127:0] out3142; 
reg [127:0] out3143; 
reg [127:0] out3144; 
reg [127:0] out3145; 
reg [127:0] out3146; 
reg [127:0] out3147; 
reg [127:0] out3148; 
reg [127:0] out3149; 
reg [127:0] out3150; 
reg [127:0] out3151; 
reg [127:0] out3152; 
reg [127:0] out3153; 
reg [127:0] out3154; 
reg [127:0] out3155; 
reg [127:0] out3156; 
reg [127:0] out3157; 
reg [127:0] out3158; 
reg [127:0] out3159; 
reg [127:0] out3160; 
reg [127:0] out3161; 
reg [127:0] out3162; 
reg [127:0] out3163; 
reg [127:0] out3164; 
reg [127:0] out3165; 
reg [127:0] out3166; 
reg [127:0] out3167; 
reg [127:0] out3168; 
reg [127:0] out3169; 
reg [127:0] out3170; 
reg [127:0] out3171; 
reg [127:0] out3172; 
reg [127:0] out3173; 
reg [127:0] out3174; 
reg [127:0] out3175; 
reg [127:0] out3176; 
reg [127:0] out3177; 
reg [127:0] out3178; 
reg [127:0] out3179; 
reg [127:0] out3180; 
reg [127:0] out3181; 
reg [127:0] out3182; 
reg [127:0] out3183; 
reg [127:0] out3184; 
reg [127:0] out3185; 
reg [127:0] out3186; 
reg [127:0] out3187; 
reg [127:0] out3188; 
reg [127:0] out3189; 
reg [127:0] out3190; 
reg [127:0] out3191; 
reg [127:0] out3192; 
reg [127:0] out3193; 
reg [127:0] out3194; 
reg [127:0] out3195; 
reg [127:0] out3196; 
reg [127:0] out3197; 
reg [127:0] out3198; 
reg [127:0] out3199; 
reg [127:0] out3200; 
reg [127:0] out3201; 
reg [127:0] out3202; 
reg [127:0] out3203; 
reg [127:0] out3204; 
reg [127:0] out3205; 
reg [127:0] out3206; 
reg [127:0] out3207; 
reg [127:0] out3208; 
reg [127:0] out3209; 
reg [127:0] out3210; 
reg [127:0] out3211; 
reg [127:0] out3212; 
reg [127:0] out3213; 
reg [127:0] out3214; 
reg [127:0] out3215; 
reg [127:0] out3216; 
reg [127:0] out3217; 
reg [127:0] out3218; 
reg [127:0] out3219; 
reg [127:0] out3220; 
reg [127:0] out3221; 
reg [127:0] out3222; 
reg [127:0] out3223; 
reg [127:0] out3224; 
reg [127:0] out3225; 
reg [127:0] out3226; 
reg [127:0] out3227; 
reg [127:0] out3228; 
reg [127:0] out3229; 
reg [127:0] out3230; 
reg [127:0] out3231; 
reg [127:0] out3232; 
reg [127:0] out3233; 
reg [127:0] out3234; 
reg [127:0] out3235; 
reg [127:0] out3236; 
reg [127:0] out3237; 
reg [127:0] out3238; 
reg [127:0] out3239; 
reg [127:0] out3240; 
reg [127:0] out3241; 
reg [127:0] out3242; 
reg [127:0] out3243; 
reg [127:0] out3244; 
reg [127:0] out3245; 
reg [127:0] out3246; 
reg [127:0] out3247; 
reg [127:0] out3248; 
reg [127:0] out3249; 
reg [127:0] out3250; 
reg [127:0] out3251; 
reg [127:0] out3252; 
reg [127:0] out3253; 
reg [127:0] out3254; 
reg [127:0] out3255; 
reg [127:0] out3256; 
reg [127:0] out3257; 
reg [127:0] out3258; 
reg [127:0] out3259; 
reg [127:0] out3260; 
reg [127:0] out3261; 
reg [127:0] out3262; 
reg [127:0] out3263; 
reg [127:0] out3264; 
reg [127:0] out3265; 
reg [127:0] out3266; 
reg [127:0] out3267; 
reg [127:0] out3268; 
reg [127:0] out3269; 
reg [127:0] out3270; 
reg [127:0] out3271; 
reg [127:0] out3272; 
reg [127:0] out3273; 
reg [127:0] out3274; 
reg [127:0] out3275; 
reg [127:0] out3276; 
reg [127:0] out3277; 
reg [127:0] out3278; 
reg [127:0] out3279; 
reg [127:0] out3280; 
reg [127:0] out3281; 
reg [127:0] out3282; 
reg [127:0] out3283; 
reg [127:0] out3284; 
reg [127:0] out3285; 
reg [127:0] out3286; 
reg [127:0] out3287; 
reg [127:0] out3288; 
reg [127:0] out3289; 
reg [127:0] out3290; 
reg [127:0] out3291; 
reg [127:0] out3292; 
reg [127:0] out3293; 
reg [127:0] out3294; 
reg [127:0] out3295; 
reg [127:0] out3296; 
reg [127:0] out3297; 
reg [127:0] out3298; 
reg [127:0] out3299; 
reg [127:0] out3300; 
reg [127:0] out3301; 
reg [127:0] out3302; 
reg [127:0] out3303; 
reg [127:0] out3304; 
reg [127:0] out3305; 
reg [127:0] out3306; 
reg [127:0] out3307; 
reg [127:0] out3308; 
reg [127:0] out3309; 
reg [127:0] out3310; 
reg [127:0] out3311; 
reg [127:0] out3312; 
reg [127:0] out3313; 
reg [127:0] out3314; 
reg [127:0] out3315; 
reg [127:0] out3316; 
reg [127:0] out3317; 
reg [127:0] out3318; 
reg [127:0] out3319; 
reg [127:0] out3320; 
reg [127:0] out3321; 
reg [127:0] out3322; 
reg [127:0] out3323; 
reg [127:0] out3324; 
reg [127:0] out3325; 
reg [127:0] out3326; 
reg [127:0] out3327; 
reg [127:0] out3328; 
reg [127:0] out3329; 
reg [127:0] out3330; 
reg [127:0] out3331; 
reg [127:0] out3332; 
reg [127:0] out3333; 
reg [127:0] out3334; 
reg [127:0] out3335; 
reg [127:0] out3336; 
reg [127:0] out3337; 
reg [127:0] out3338; 
reg [127:0] out3339; 
reg [127:0] out3340; 
reg [127:0] out3341; 
reg [127:0] out3342; 
reg [127:0] out3343; 
reg [127:0] out3344; 
reg [127:0] out3345; 
reg [127:0] out3346; 
reg [127:0] out3347; 
reg [127:0] out3348; 
reg [127:0] out3349; 
reg [127:0] out3350; 
reg [127:0] out3351; 
reg [127:0] out3352; 
reg [127:0] out3353; 
reg [127:0] out3354; 
reg [127:0] out3355; 
reg [127:0] out3356; 
reg [127:0] out3357; 
reg [127:0] out3358; 
reg [127:0] out3359; 
reg [127:0] out3360; 
reg [127:0] out3361; 
reg [127:0] out3362; 
reg [127:0] out3363; 
reg [127:0] out3364; 
reg [127:0] out3365; 
reg [127:0] out3366; 
reg [127:0] out3367; 
reg [127:0] out3368; 
reg [127:0] out3369; 
reg [127:0] out3370; 
reg [127:0] out3371; 
reg [127:0] out3372; 
reg [127:0] out3373; 
reg [127:0] out3374; 
reg [127:0] out3375; 
reg [127:0] out3376; 
reg [127:0] out3377; 
reg [127:0] out3378; 
reg [127:0] out3379; 
reg [127:0] out3380; 
reg [127:0] out3381; 
reg [127:0] out3382; 
reg [127:0] out3383; 
reg [127:0] out3384; 
reg [127:0] out3385; 
reg [127:0] out3386; 
reg [127:0] out3387; 
reg [127:0] out3388; 
reg [127:0] out3389; 
reg [127:0] out3390; 
reg [127:0] out3391; 
reg [127:0] out3392; 
reg [127:0] out3393; 
reg [127:0] out3394; 
reg [127:0] out3395; 
reg [127:0] out3396; 
reg [127:0] out3397; 
reg [127:0] out3398; 
reg [127:0] out3399; 
reg [127:0] out3400; 
reg [127:0] out3401; 
reg [127:0] out3402; 
reg [127:0] out3403; 
reg [127:0] out3404; 
reg [127:0] out3405; 
reg [127:0] out3406; 
reg [127:0] out3407; 
reg [127:0] out3408; 
reg [127:0] out3409; 
reg [127:0] out3410; 
reg [127:0] out3411; 
reg [127:0] out3412; 
reg [127:0] out3413; 
reg [127:0] out3414; 
reg [127:0] out3415; 
reg [127:0] out3416; 
reg [127:0] out3417; 
reg [127:0] out3418; 
reg [127:0] out3419; 
reg [127:0] out3420; 
reg [127:0] out3421; 
reg [127:0] out3422; 
reg [127:0] out3423; 
reg [127:0] out3424; 
reg [127:0] out3425; 
reg [127:0] out3426; 
reg [127:0] out3427; 
reg [127:0] out3428; 
reg [127:0] out3429; 
reg [127:0] out3430; 
reg [127:0] out3431; 
reg [127:0] out3432; 
reg [127:0] out3433; 
reg [127:0] out3434; 
reg [127:0] out3435; 
reg [127:0] out3436; 
reg [127:0] out3437; 
reg [127:0] out3438; 
reg [127:0] out3439; 
reg [127:0] out3440; 
reg [127:0] out3441; 
reg [127:0] out3442; 
reg [127:0] out3443; 
reg [127:0] out3444; 
reg [127:0] out3445; 
reg [127:0] out3446; 
reg [127:0] out3447; 
reg [127:0] out3448; 
reg [127:0] out3449; 
reg [127:0] out3450; 
reg [127:0] out3451; 
reg [127:0] out3452; 
reg [127:0] out3453; 
reg [127:0] out3454; 
reg [127:0] out3455; 
reg [127:0] out3456; 
reg [127:0] out3457; 
reg [127:0] out3458; 
reg [127:0] out3459; 
reg [127:0] out3460; 
reg [127:0] out3461; 
reg [127:0] out3462; 
reg [127:0] out3463; 
reg [127:0] out3464; 
reg [127:0] out3465; 
reg [127:0] out3466; 
reg [127:0] out3467; 
reg [127:0] out3468; 
reg [127:0] out3469; 
reg [127:0] out3470; 
reg [127:0] out3471; 
reg [127:0] out3472; 
reg [127:0] out3473; 
reg [127:0] out3474; 
reg [127:0] out3475; 
reg [127:0] out3476; 
reg [127:0] out3477; 
reg [127:0] out3478; 
reg [127:0] out3479; 
reg [127:0] out3480; 
reg [127:0] out3481; 
reg [127:0] out3482; 
reg [127:0] out3483; 
reg [127:0] out3484; 
reg [127:0] out3485; 
reg [127:0] out3486; 
reg [127:0] out3487; 
reg [127:0] out3488; 
reg [127:0] out3489; 
reg [127:0] out3490; 
reg [127:0] out3491; 
reg [127:0] out3492; 
reg [127:0] out3493; 
reg [127:0] out3494; 
reg [127:0] out3495; 
reg [127:0] out3496; 
reg [127:0] out3497; 
reg [127:0] out3498; 
reg [127:0] out3499; 
reg [127:0] out3500; 
reg [127:0] out3501; 
reg [127:0] out3502; 
reg [127:0] out3503; 
reg [127:0] out3504; 
reg [127:0] out3505; 
reg [127:0] out3506; 
reg [127:0] out3507; 
reg [127:0] out3508; 
reg [127:0] out3509; 
reg [127:0] out3510; 
reg [127:0] out3511; 
reg [127:0] out3512; 
reg [127:0] out3513; 
reg [127:0] out3514; 
reg [127:0] out3515; 
reg [127:0] out3516; 
reg [127:0] out3517; 
reg [127:0] out3518; 
reg [127:0] out3519; 
reg [127:0] out3520; 
reg [127:0] out3521; 
reg [127:0] out3522; 
reg [127:0] out3523; 
reg [127:0] out3524; 
reg [127:0] out3525; 
reg [127:0] out3526; 
reg [127:0] out3527; 
reg [127:0] out3528; 
reg [127:0] out3529; 
reg [127:0] out3530; 
reg [127:0] out3531; 
reg [127:0] out3532; 
reg [127:0] out3533; 
reg [127:0] out3534; 
reg [127:0] out3535; 
reg [127:0] out3536; 
reg [127:0] out3537; 
reg [127:0] out3538; 
reg [127:0] out3539; 
reg [127:0] out3540; 
reg [127:0] out3541; 
reg [127:0] out3542; 
reg [127:0] out3543; 
reg [127:0] out3544; 
reg [127:0] out3545; 
reg [127:0] out3546; 
reg [127:0] out3547; 
reg [127:0] out3548; 
reg [127:0] out3549; 
reg [127:0] out3550; 
reg [127:0] out3551; 
reg [127:0] out3552; 
reg [127:0] out3553; 
reg [127:0] out3554; 
reg [127:0] out3555; 
reg [127:0] out3556; 
reg [127:0] out3557; 
reg [127:0] out3558; 
reg [127:0] out3559; 
reg [127:0] out3560; 
reg [127:0] out3561; 
reg [127:0] out3562; 
reg [127:0] out3563; 
reg [127:0] out3564; 
reg [127:0] out3565; 
reg [127:0] out3566; 
reg [127:0] out3567; 
reg [127:0] out3568; 
reg [127:0] out3569; 
reg [127:0] out3570; 
reg [127:0] out3571; 
reg [127:0] out3572; 
reg [127:0] out3573; 
reg [127:0] out3574; 
reg [127:0] out3575; 
reg [127:0] out3576; 
reg [127:0] out3577; 
reg [127:0] out3578; 
reg [127:0] out3579; 
reg [127:0] out3580; 
reg [127:0] out3581; 
reg [127:0] out3582; 
reg [127:0] out3583; 
reg [127:0] out3584; 
reg [127:0] out3585; 
reg [127:0] out3586; 
reg [127:0] out3587; 
reg [127:0] out3588; 
reg [127:0] out3589; 
reg [127:0] out3590; 
reg [127:0] out3591; 
reg [127:0] out3592; 
reg [127:0] out3593; 
reg [127:0] out3594; 
reg [127:0] out3595; 
reg [127:0] out3596; 
reg [127:0] out3597; 
reg [127:0] out3598; 
reg [127:0] out3599; 
reg [127:0] out3600; 
reg [127:0] out3601; 
reg [127:0] out3602; 
reg [127:0] out3603; 
reg [127:0] out3604; 
reg [127:0] out3605; 
reg [127:0] out3606; 
reg [127:0] out3607; 
reg [127:0] out3608; 
reg [127:0] out3609; 
reg [127:0] out3610; 
reg [127:0] out3611; 
reg [127:0] out3612; 
reg [127:0] out3613; 
reg [127:0] out3614; 
reg [127:0] out3615; 
reg [127:0] out3616; 
reg [127:0] out3617; 
reg [127:0] out3618; 
reg [127:0] out3619; 
reg [127:0] out3620; 
reg [127:0] out3621; 
reg [127:0] out3622; 
reg [127:0] out3623; 
reg [127:0] out3624; 
reg [127:0] out3625; 
reg [127:0] out3626; 
reg [127:0] out3627; 
reg [127:0] out3628; 
reg [127:0] out3629; 
reg [127:0] out3630; 
reg [127:0] out3631; 
reg [127:0] out3632; 
reg [127:0] out3633; 
reg [127:0] out3634; 
reg [127:0] out3635; 
reg [127:0] out3636; 
reg [127:0] out3637; 
reg [127:0] out3638; 
reg [127:0] out3639; 
reg [127:0] out3640; 
reg [127:0] out3641; 
reg [127:0] out3642; 
reg [127:0] out3643; 
reg [127:0] out3644; 
reg [127:0] out3645; 
reg [127:0] out3646; 
reg [127:0] out3647; 
reg [127:0] out3648; 
reg [127:0] out3649; 
reg [127:0] out3650; 
reg [127:0] out3651; 
reg [127:0] out3652; 
reg [127:0] out3653; 
reg [127:0] out3654; 
reg [127:0] out3655; 
reg [127:0] out3656; 
reg [127:0] out3657; 
reg [127:0] out3658; 
reg [127:0] out3659; 
reg [127:0] out3660; 
reg [127:0] out3661; 
reg [127:0] out3662; 
reg [127:0] out3663; 
reg [127:0] out3664; 
reg [127:0] out3665; 
reg [127:0] out3666; 
reg [127:0] out3667; 
reg [127:0] out3668; 
reg [127:0] out3669; 
reg [127:0] out3670; 
reg [127:0] out3671; 
reg [127:0] out3672; 
reg [127:0] out3673; 
reg [127:0] out3674; 
reg [127:0] out3675; 
reg [127:0] out3676; 
reg [127:0] out3677; 
reg [127:0] out3678; 
reg [127:0] out3679; 
reg [127:0] out3680; 
reg [127:0] out3681; 
reg [127:0] out3682; 
reg [127:0] out3683; 
reg [127:0] out3684; 
reg [127:0] out3685; 
reg [127:0] out3686; 
reg [127:0] out3687; 
reg [127:0] out3688; 
reg [127:0] out3689; 
reg [127:0] out3690; 
reg [127:0] out3691; 
reg [127:0] out3692; 
reg [127:0] out3693; 
reg [127:0] out3694; 
reg [127:0] out3695; 
reg [127:0] out3696; 
reg [127:0] out3697; 
reg [127:0] out3698; 
reg [127:0] out3699; 
reg [127:0] out3700; 
reg [127:0] out3701; 
reg [127:0] out3702; 
reg [127:0] out3703; 
reg [127:0] out3704; 
reg [127:0] out3705; 
reg [127:0] out3706; 
reg [127:0] out3707; 
reg [127:0] out3708; 
reg [127:0] out3709; 
reg [127:0] out3710; 
reg [127:0] out3711; 
reg [127:0] out3712; 
reg [127:0] out3713; 
reg [127:0] out3714; 
reg [127:0] out3715; 
reg [127:0] out3716; 
reg [127:0] out3717; 
reg [127:0] out3718; 
reg [127:0] out3719; 
reg [127:0] out3720; 
reg [127:0] out3721; 
reg [127:0] out3722; 
reg [127:0] out3723; 
reg [127:0] out3724; 
reg [127:0] out3725; 
reg [127:0] out3726; 
reg [127:0] out3727; 
reg [127:0] out3728; 
reg [127:0] out3729; 
reg [127:0] out3730; 
reg [127:0] out3731; 
reg [127:0] out3732; 
reg [127:0] out3733; 
reg [127:0] out3734; 
reg [127:0] out3735; 
reg [127:0] out3736; 
reg [127:0] out3737; 
reg [127:0] out3738; 
reg [127:0] out3739; 
reg [127:0] out3740; 
reg [127:0] out3741; 
reg [127:0] out3742; 
reg [127:0] out3743; 
reg [127:0] out3744; 
reg [127:0] out3745; 
reg [127:0] out3746; 
reg [127:0] out3747; 
reg [127:0] out3748; 
reg [127:0] out3749; 
reg [127:0] out3750; 
reg [127:0] out3751; 
reg [127:0] out3752; 
reg [127:0] out3753; 
reg [127:0] out3754; 
reg [127:0] out3755; 
reg [127:0] out3756; 
reg [127:0] out3757; 
reg [127:0] out3758; 
reg [127:0] out3759; 
reg [127:0] out3760; 
reg [127:0] out3761; 
reg [127:0] out3762; 
reg [127:0] out3763; 
reg [127:0] out3764; 
reg [127:0] out3765; 
reg [127:0] out3766; 
reg [127:0] out3767; 
reg [127:0] out3768; 
reg [127:0] out3769; 
reg [127:0] out3770; 
reg [127:0] out3771; 
reg [127:0] out3772; 
reg [127:0] out3773; 
reg [127:0] out3774; 
reg [127:0] out3775; 
reg [127:0] out3776; 
reg [127:0] out3777; 
reg [127:0] out3778; 
reg [127:0] out3779; 
reg [127:0] out3780; 
reg [127:0] out3781; 
reg [127:0] out3782; 
reg [127:0] out3783; 
reg [127:0] out3784; 
reg [127:0] out3785; 
reg [127:0] out3786; 
reg [127:0] out3787; 
reg [127:0] out3788; 
reg [127:0] out3789; 
reg [127:0] out3790; 
reg [127:0] out3791; 
reg [127:0] out3792; 
reg [127:0] out3793; 
reg [127:0] out3794; 
reg [127:0] out3795; 
reg [127:0] out3796; 
reg [127:0] out3797; 
reg [127:0] out3798; 
reg [127:0] out3799; 
reg [127:0] out3800; 
reg [127:0] out3801; 
reg [127:0] out3802; 
reg [127:0] out3803; 
reg [127:0] out3804; 
reg [127:0] out3805; 
reg [127:0] out3806; 
reg [127:0] out3807; 
reg [127:0] out3808; 
reg [127:0] out3809; 
reg [127:0] out3810; 
reg [127:0] out3811; 
reg [127:0] out3812; 
reg [127:0] out3813; 
reg [127:0] out3814; 
reg [127:0] out3815; 
reg [127:0] out3816; 
reg [127:0] out3817; 
reg [127:0] out3818; 
reg [127:0] out3819; 
reg [127:0] out3820; 
reg [127:0] out3821; 
reg [127:0] out3822; 
reg [127:0] out3823; 
reg [127:0] out3824; 
reg [127:0] out3825; 
reg [127:0] out3826; 
reg [127:0] out3827; 
reg [127:0] out3828; 
reg [127:0] out3829; 
reg [127:0] out3830; 
reg [127:0] out3831; 
reg [127:0] out3832; 
reg [127:0] out3833; 
reg [127:0] out3834; 
reg [127:0] out3835; 
reg [127:0] out3836; 
reg [127:0] out3837; 
reg [127:0] out3838; 
reg [127:0] out3839; 
reg [127:0] out3840; 
reg [127:0] out3841; 
reg [127:0] out3842; 
reg [127:0] out3843; 
reg [127:0] out3844; 
reg [127:0] out3845; 
reg [127:0] out3846; 
reg [127:0] out3847; 
reg [127:0] out3848; 
reg [127:0] out3849; 
reg [127:0] out3850; 
reg [127:0] out3851; 
reg [127:0] out3852; 
reg [127:0] out3853; 
reg [127:0] out3854; 
reg [127:0] out3855; 
reg [127:0] out3856; 
reg [127:0] out3857; 
reg [127:0] out3858; 
reg [127:0] out3859; 
reg [127:0] out3860; 
reg [127:0] out3861; 
reg [127:0] out3862; 
reg [127:0] out3863; 
reg [127:0] out3864; 
reg [127:0] out3865; 
reg [127:0] out3866; 
reg [127:0] out3867; 
reg [127:0] out3868; 
reg [127:0] out3869; 
reg [127:0] out3870; 
reg [127:0] out3871; 
reg [127:0] out3872; 
reg [127:0] out3873; 
reg [127:0] out3874; 
reg [127:0] out3875; 
reg [127:0] out3876; 
reg [127:0] out3877; 
reg [127:0] out3878; 
reg [127:0] out3879; 
reg [127:0] out3880; 
reg [127:0] out3881; 
reg [127:0] out3882; 
reg [127:0] out3883; 
reg [127:0] out3884; 
reg [127:0] out3885; 
reg [127:0] out3886; 
reg [127:0] out3887; 
reg [127:0] out3888; 
reg [127:0] out3889; 
reg [127:0] out3890; 
reg [127:0] out3891; 
reg [127:0] out3892; 
reg [127:0] out3893; 
reg [127:0] out3894; 
reg [127:0] out3895; 
reg [127:0] out3896; 
reg [127:0] out3897; 
reg [127:0] out3898; 
reg [127:0] out3899; 
reg [127:0] out3900; 
reg [127:0] out3901; 
reg [127:0] out3902; 
reg [127:0] out3903; 
reg [127:0] out3904; 
reg [127:0] out3905; 
reg [127:0] out3906; 
reg [127:0] out3907; 
reg [127:0] out3908; 
reg [127:0] out3909; 
reg [127:0] out3910; 
reg [127:0] out3911; 
reg [127:0] out3912; 
reg [127:0] out3913; 
reg [127:0] out3914; 
reg [127:0] out3915; 
reg [127:0] out3916; 
reg [127:0] out3917; 
reg [127:0] out3918; 
reg [127:0] out3919; 
reg [127:0] out3920; 
reg [127:0] out3921; 
reg [127:0] out3922; 
reg [127:0] out3923; 
reg [127:0] out3924; 
reg [127:0] out3925; 
reg [127:0] out3926; 
reg [127:0] out3927; 
reg [127:0] out3928; 
reg [127:0] out3929; 
reg [127:0] out3930; 
reg [127:0] out3931; 
reg [127:0] out3932; 
reg [127:0] out3933; 
reg [127:0] out3934; 
reg [127:0] out3935; 
reg [127:0] out3936; 
reg [127:0] out3937; 
reg [127:0] out3938; 
reg [127:0] out3939; 
reg [127:0] out3940; 
reg [127:0] out3941; 
reg [127:0] out3942; 
reg [127:0] out3943; 
reg [127:0] out3944; 
reg [127:0] out3945; 
reg [127:0] out3946; 
reg [127:0] out3947; 
reg [127:0] out3948; 
reg [127:0] out3949; 
reg [127:0] out3950; 
reg [127:0] out3951; 
reg [127:0] out3952; 
reg [127:0] out3953; 
reg [127:0] out3954; 
reg [127:0] out3955; 
reg [127:0] out3956; 
reg [127:0] out3957; 
reg [127:0] out3958; 
reg [127:0] out3959; 
reg [127:0] out3960; 
reg [127:0] out3961; 
reg [127:0] out3962; 
reg [127:0] out3963; 
reg [127:0] out3964; 
reg [127:0] out3965; 
reg [127:0] out3966; 
reg [127:0] out3967; 
reg [127:0] out3968; 
reg [127:0] out3969; 
reg [127:0] out3970; 
reg [127:0] out3971; 
reg [127:0] out3972; 
reg [127:0] out3973; 
reg [127:0] out3974; 
reg [127:0] out3975; 
reg [127:0] out3976; 
reg [127:0] out3977; 
reg [127:0] out3978; 
reg [127:0] out3979; 
reg [127:0] out3980; 
reg [127:0] out3981; 
reg [127:0] out3982; 
reg [127:0] out3983; 
reg [127:0] out3984; 
reg [127:0] out3985; 
reg [127:0] out3986; 
reg [127:0] out3987; 
reg [127:0] out3988; 
reg [127:0] out3989; 
reg [127:0] out3990; 
reg [127:0] out3991; 
reg [127:0] out3992; 
reg [127:0] out3993; 
reg [127:0] out3994; 
reg [127:0] out3995; 
reg [127:0] out3996; 
reg [127:0] out3997; 
reg [127:0] out3998; 
reg [127:0] out3999; 
reg [127:0] out4000; 
reg [127:0] out4001; 
reg [127:0] out4002; 
reg [127:0] out4003; 
reg [127:0] out4004; 
reg [127:0] out4005; 
reg [127:0] out4006; 
reg [127:0] out4007; 
reg [127:0] out4008; 
reg [127:0] out4009; 
reg [127:0] out4010; 
reg [127:0] out4011; 
reg [127:0] out4012; 
reg [127:0] out4013; 
reg [127:0] out4014; 
reg [127:0] out4015; 
reg [127:0] out4016; 
reg [127:0] out4017; 
reg [127:0] out4018; 
reg [127:0] out4019; 
reg [127:0] out4020; 
reg [127:0] out4021; 
reg [127:0] out4022; 
reg [127:0] out4023; 
reg [127:0] out4024; 
reg [127:0] out4025; 
reg [127:0] out4026; 
reg [127:0] out4027; 
reg [127:0] out4028; 
reg [127:0] out4029; 
reg [127:0] out4030; 
reg [127:0] out4031; 
reg [127:0] out4032; 
reg [127:0] out4033; 
reg [127:0] out4034; 
reg [127:0] out4035; 
reg [127:0] out4036; 
reg [127:0] out4037; 
reg [127:0] out4038; 
reg [127:0] out4039; 
reg [127:0] out4040; 
reg [127:0] out4041; 
reg [127:0] out4042; 
reg [127:0] out4043; 
reg [127:0] out4044; 
reg [127:0] out4045; 
reg [127:0] out4046; 
reg [127:0] out4047; 
reg [127:0] out4048; 
reg [127:0] out4049; 
reg [127:0] out4050; 
reg [127:0] out4051; 
reg [127:0] out4052; 
reg [127:0] out4053; 
reg [127:0] out4054; 
reg [127:0] out4055; 
reg [127:0] out4056; 
reg [127:0] out4057; 
reg [127:0] out4058; 
reg [127:0] out4059; 
reg [127:0] out4060; 
reg [127:0] out4061; 
reg [127:0] out4062; 
reg [127:0] out4063; 
reg [127:0] out4064; 
reg [127:0] out4065; 
reg [127:0] out4066; 
reg [127:0] out4067; 
reg [127:0] out4068; 
reg [127:0] out4069; 
reg [127:0] out4070; 
reg [127:0] out4071; 
reg [127:0] out4072; 
reg [127:0] out4073; 
reg [127:0] out4074; 
reg [127:0] out4075; 
reg [127:0] out4076; 
reg [127:0] out4077; 
reg [127:0] out4078; 
reg [127:0] out4079; 
reg [127:0] out4080; 
reg [127:0] out4081; 
reg [127:0] out4082; 
reg [127:0] out4083; 
reg [127:0] out4084; 
reg [127:0] out4085; 
reg [127:0] out4086; 
reg [127:0] out4087; 
reg [127:0] out4088; 
reg [127:0] out4089; 
reg [127:0] out4090; 
reg [127:0] out4091; 
reg [127:0] out4092; 
reg [127:0] out4093; 
reg [127:0] out4094; 
reg [127:0] out4095; 
reg [127:0] out4096; 
reg [127:0] out4097; 
reg [127:0] out4098; 
reg [127:0] out4099; 
reg [127:0] out4100; 
reg [127:0] out4101; 
reg [127:0] out4102; 
reg [127:0] out4103; 
reg [127:0] out4104; 
reg [127:0] out4105; 
reg [127:0] out4106; 
reg [127:0] out4107; 
reg [127:0] out4108; 
reg [127:0] out4109; 
reg [127:0] out4110; 
reg [127:0] out4111; 
reg [127:0] out4112; 
reg [127:0] out4113; 
reg [127:0] out4114; 
reg [127:0] out4115; 
reg [127:0] out4116; 
reg [127:0] out4117; 
reg [127:0] out4118; 
reg [127:0] out4119; 
reg [127:0] out4120; 
reg [127:0] out4121; 
reg [127:0] out4122; 
reg [127:0] out4123; 
reg [127:0] out4124; 
reg [127:0] out4125; 
reg [127:0] out4126; 
reg [127:0] out4127; 
reg [127:0] out4128; 
reg [127:0] out4129; 
reg [127:0] out4130; 
reg [127:0] out4131; 
reg [127:0] out4132; 
reg [127:0] out4133; 
reg [127:0] out4134; 
reg [127:0] out4135; 
reg [127:0] out4136; 
reg [127:0] out4137; 
reg [127:0] out4138; 
reg [127:0] out4139; 
reg [127:0] out4140; 
reg [127:0] out4141; 
reg [127:0] out4142; 
reg [127:0] out4143; 
reg [127:0] out4144; 
reg [127:0] out4145; 
reg [127:0] out4146; 
reg [127:0] out4147; 
reg [127:0] out4148; 
reg [127:0] out4149; 
reg [127:0] out4150; 
reg [127:0] out4151; 
reg [127:0] out4152; 
reg [127:0] out4153; 
reg [127:0] out4154; 
reg [127:0] out4155; 
reg [127:0] out4156; 
reg [127:0] out4157; 
reg [127:0] out4158; 
reg [127:0] out4159; 
reg [127:0] out4160; 
reg [127:0] out4161; 
reg [127:0] out4162; 
reg [127:0] out4163; 
reg [127:0] out4164; 
reg [127:0] out4165; 
reg [127:0] out4166; 
reg [127:0] out4167; 
reg [127:0] out4168; 
reg [127:0] out4169; 
reg [127:0] out4170; 
reg [127:0] out4171; 
reg [127:0] out4172; 
reg [127:0] out4173; 
reg [127:0] out4174; 
reg [127:0] out4175; 
reg [127:0] out4176; 
reg [127:0] out4177; 
reg [127:0] out4178; 
reg [127:0] out4179; 
reg [127:0] out4180; 
reg [127:0] out4181; 
reg [127:0] out4182; 
reg [127:0] out4183; 
reg [127:0] out4184; 
reg [127:0] out4185; 
reg [127:0] out4186; 
reg [127:0] out4187; 
reg [127:0] out4188; 
reg [127:0] out4189; 
reg [127:0] out4190; 
reg [127:0] out4191; 
reg [127:0] out4192; 
reg [127:0] out4193; 
reg [127:0] out4194; 
reg [127:0] out4195; 
reg [127:0] out4196; 
reg [127:0] out4197; 
reg [127:0] out4198; 
reg [127:0] out4199; 
reg [127:0] out4200; 
reg [127:0] out4201; 
reg [127:0] out4202; 
reg [127:0] out4203; 
reg [127:0] out4204; 
reg [127:0] out4205; 
reg [127:0] out4206; 
reg [127:0] out4207; 
reg [127:0] out4208; 
reg [127:0] out4209; 
reg [127:0] out4210; 
reg [127:0] out4211; 
reg [127:0] out4212; 
reg [127:0] out4213; 
reg [127:0] out4214; 
reg [127:0] out4215; 
reg [127:0] out4216; 
reg [127:0] out4217; 
reg [127:0] out4218; 
reg [127:0] out4219; 
reg [127:0] out4220; 
reg [127:0] out4221; 
reg [127:0] out4222; 
reg [127:0] out4223; 
reg [127:0] out4224; 
reg [127:0] out4225; 
reg [127:0] out4226; 
reg [127:0] out4227; 
reg [127:0] out4228; 
reg [127:0] out4229; 
reg [127:0] out4230; 
reg [127:0] out4231; 
reg [127:0] out4232; 
reg [127:0] out4233; 
reg [127:0] out4234; 
reg [127:0] out4235; 
reg [127:0] out4236; 
reg [127:0] out4237; 
reg [127:0] out4238; 
reg [127:0] out4239; 
reg [127:0] out4240; 
reg [127:0] out4241; 
reg [127:0] out4242; 
reg [127:0] out4243; 
reg [127:0] out4244; 
reg [127:0] out4245; 
reg [127:0] out4246; 
reg [127:0] out4247; 
reg [127:0] out4248; 
reg [127:0] out4249; 
reg [127:0] out4250; 
reg [127:0] out4251; 
reg [127:0] out4252; 
reg [127:0] out4253; 
reg [127:0] out4254; 
reg [127:0] out4255; 
reg [127:0] out4256; 
reg [127:0] out4257; 
reg [127:0] out4258; 
reg [127:0] out4259; 
reg [127:0] out4260; 
reg [127:0] out4261; 
reg [127:0] out4262; 
reg [127:0] out4263; 
reg [127:0] out4264; 
reg [127:0] out4265; 
reg [127:0] out4266; 
reg [127:0] out4267; 
reg [127:0] out4268; 
reg [127:0] out4269; 
reg [127:0] out4270; 
reg [127:0] out4271; 
reg [127:0] out4272; 
reg [127:0] out4273; 
reg [127:0] out4274; 
reg [127:0] out4275; 
reg [127:0] out4276; 
reg [127:0] out4277; 
reg [127:0] out4278; 
reg [127:0] out4279; 
reg [127:0] out4280; 
reg [127:0] out4281; 
reg [127:0] out4282; 
reg [127:0] out4283; 
reg [127:0] out4284; 
reg [127:0] out4285; 
reg [127:0] out4286; 
reg [127:0] out4287; 
reg [127:0] out4288; 
reg [127:0] out4289; 
reg [127:0] out4290; 
reg [127:0] out4291; 
reg [127:0] out4292; 
reg [127:0] out4293; 
reg [127:0] out4294; 
reg [127:0] out4295; 
reg [127:0] out4296; 
reg [127:0] out4297; 
reg [127:0] out4298; 
reg [127:0] out4299; 
reg [127:0] out4300; 
reg [127:0] out4301; 
reg [127:0] out4302; 
reg [127:0] out4303; 
reg [127:0] out4304; 
reg [127:0] out4305; 
reg [127:0] out4306; 
reg [127:0] out4307; 
reg [127:0] out4308; 
reg [127:0] out4309; 
reg [127:0] out4310; 
reg [127:0] out4311; 
reg [127:0] out4312; 
reg [127:0] out4313; 
reg [127:0] out4314; 
reg [127:0] out4315; 
reg [127:0] out4316; 
reg [127:0] out4317; 
reg [127:0] out4318; 
reg [127:0] out4319; 
reg [127:0] out4320; 
reg [127:0] out4321; 
reg [127:0] out4322; 
reg [127:0] out4323; 
reg [127:0] out4324; 
reg [127:0] out4325; 
reg [127:0] out4326; 
reg [127:0] out4327; 
reg [127:0] out4328; 
reg [127:0] out4329; 
reg [127:0] out4330; 
reg [127:0] out4331; 
reg [127:0] out4332; 
reg [127:0] out4333; 
reg [127:0] out4334; 
reg [127:0] out4335; 
reg [127:0] out4336; 
reg [127:0] out4337; 
reg [127:0] out4338; 
reg [127:0] out4339; 
reg [127:0] out4340; 
top uut ( 
.clk(clk), 
.rst(rst), 
.state(state), 
.key(key), 
.out(out), 
.Antena(Antena) 
); 
initial begin 
f = $fopen("data_0.000_00_2.csv","a"); 
clk = 0; 
state = 0; 
key = 0; 
bit_err = 128'b0; 
@ (negedge clk); 
#20;
rst = 1;
$fwrite(f,"%b, %b, %b, %b\n",state, out1, out, Antena); 
@ (negedge clk); 
#20;
rst = 0;
$fwrite(f,"%b, %b, %b, %b\n",state, out1, out, Antena); 		
#60; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111110001010100111001001000011000001110010000011001101001101100001110011001010110100001011100011011001011000101110010110000; 
out1 = 128'b00010000100111011000010100001101100111110010000101111001011000101000011111011100011010001010001101000101010110100000110101000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110100101101110001100100110100111101010000110011111010000010110100111100001101100111000110100010111001110000111110011110010; 
out2 = 128'b11101001110100000101100111101001000101100110110001001111001101011010000100110101011110100101000010001010100011111100111010010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011111111111101010100101000011001011001100000101010000100011101111011000111110110011010111000111111100011000000110011000010; 
out3 = 128'b00100100001001010011110001001111000111110101001101000100101011000011011011100000001101011100111111100100110001101010111111101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001001011100110111001001101011101000110100000111011101111110000001101101011011010101110100100010100110101100001101101111110000; 
out4 = 128'b11011101011111001111011000010000010100010011011011111110011101001110101000100110100101100000000101101110010111001110000111101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101111011110010001111010011010011101010010100000000101011110011000000110011000100001100111110101101110001111100110010000100; 
out5 = 128'b11010101111111010011100101110000111100000100010101010001000010100000100010101010111100010110010011100100111011011011111010101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out5[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out5, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101101101110100110011110100111110100000001010110010110000100010100000110001001011000101010001001110001001101000001111100101110; 
out6 = 128'b00011001010101011111011111110011011010001010110000011001010001001110100011100100100011001111001111001000000101010001010010001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out6[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out6, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111111101110101011001001101010011101101001000001011110110101000010001110000011011101100100001011010101011100110100111100010; 
out7 = 128'b01110111100010011100000100000001111010000111100011101101011100000001000010100011000011111001100000111000000111000000010001111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out7[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out7, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100011100100110101100001111001110010000100110001010000110000110111010110010111011100101101100000001000011001111010100110010; 
out8 = 128'b11001001011100010011111000111101110010001010110100001101011000001010010100101111001110100111000100001011001100100001001101010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out8[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out8, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010100000111011001011110100100001000000001001110001011101010101001001011110000000100101110101000011111110010110101110100010; 
out9 = 128'b11110101001100111111111000110101101111000000001101110011111111101111001100010111011100010011010111001111011001110110110000010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out9[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out9, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110100100011110000000001010011011000010010111010111111010000100011010111111111100000100111100101010110000010011011011000100; 
out10 = 128'b10001100000100110100000100011111111000100000101111111111001111001011110011111110011011010000101010100001111110010101001110000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out10[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out10, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100001101110110001110101100000100100001111000110000110111111101101111000110110011011111001100000001111011101010011010010001; 
out11 = 128'b00110011100000001100000101011101001010010011101100001101001010101010011010010001000001100010101111001010101011010100111101001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out11[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out11, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011011011111001011101011011101010111000101100111001110111011001110011111011001101000101110000101100100010001111100011010101; 
out12 = 128'b00110111100010101101111100110000001001100011001011101101101110001001010000000011100010010101010010000011011101101111010111011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out12[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out12, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110001111000100001000110010001011101011100100000010000111110101001101110011010000101101110111010111101000101001101010111001; 
out13 = 128'b01110110100000100000110001110101100111111111011100100011011100000100010001111110110001100011000101001101101110010110010101110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out13[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out13, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000101101100101001011010110111001111111110001100011100110011001011110110111111101111001101110011010101111010100010001010111; 
out14 = 128'b10010101000111101001000110001000100101001100111101010100000100110001111000110010011101010101110010111001111100100010101101111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out14[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out14, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111111000000110101101101100111011000101001110110011011010100101011001011101100110100010111011011110001111001000110100011001; 
out15 = 128'b01100101101010101001100011010110000100101101001110011011010100110011101111011100101011001011110000001001001101100001011100011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out15[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out15, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100011001011110000000000001101100110111111110100110010010111100111100011001010010100100001100000001100101000101010111100011; 
out16 = 128'b10010110101011110110010100111111001110010100111001100000110100000111001010100101111000000001101001101111101111101111010110010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out16[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out16, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010000111111011000100010111010011101011101100001110011000010000110011100111011010011010001101110101101000001111110101011001; 
out17 = 128'b10101001001010101110011101100010010000000000111111101001100010010001110000000110101011011000100011001100101110010011110101110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out17[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out17, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100110110100101111111001101000011110101001001100100011110001101110100100010000110010010111100010001010010011101011010101001; 
out18 = 128'b10001011010001010000101100001001000011101110011111101001010000101101111011001100011011111001101110100000111011101101000010011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out18[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out18, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011100100101110101001101011001111000000110100010000101010011100000010110001101100010111110001111110111100011110111100001110; 
out19 = 128'b01001101000110101101110110011111010100000010111100010100110000010010010110101000000110100011110111100010001010001100110111010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out19[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out19, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110110100100111100110000110001001001011101110101101011000010011100100111110011111001011011111100011101101111111101000100101; 
out20 = 128'b00100100000101100001111011100100111000000001001011011100000101111000110011101101110100111010100010000111001110101110110000101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out20[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out20, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000000000000101110000001100101101011100010001110000100011000100001000001110110011111101111110111000010000011011001010110111; 
out21 = 128'b11010100000001100110001111101001101110001011101000110100110001100011100111100101011101100000010000011000101010010111010000111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out21[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out21, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110001101110110000011101010010011111010000001101110010111011111101001110111011111101100010101000101111010000000111000100111; 
out22 = 128'b11110100001110001011010110110001111001101101000101010010010010101100110000011010110111101110101111101101010011111110100000011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out22[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out22, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100101111101000100101110111100000010010000100111000111010110110001100011111110010010111010011001000011010001110101010111010; 
out23 = 128'b11010101011110010100011011011111000100110001101100110010100111000110001011010101100011010111001010001110011001100010100001101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out23[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out23, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010110000001100000011101000001111101111111000010101101111100111001100111101101111000101010111011111111110101111000111011000; 
out24 = 128'b00111000110010101100010110001111010110010011010100010100011010001011111110111111100010110101000001010000011000100001001111001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out24[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out24, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111011000100010000001000110101111010011010011011101001000100000011110111100101100011001001110011011000000111010000110111010; 
out25 = 128'b10011001110010001111000100010000001001110001100100110100110101000111100000110011010010110111011110100110000001001001011110010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out25[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out25, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010011111110100101000110001101111110100100111100101110000000111110010110000001101011010101010000111001111011000000011101101000; 
out26 = 128'b10011110101111100001010110100110010111110111110100101001100100010011001100010110010100101100001000111000100001001010001111011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out26[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out26, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001000101000011001101000110000001111011111101110011010100101101100111001100100110100101101111111011011110100010100000110111111; 
out27 = 128'b11000110111101001000010011010100100000101101110110111100000001101000111111000101110011101101010110001101001010101000101111000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out27[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out27, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000010010011110000010111101111010110110100001111110111101001000001111010101101011101010011101010110100111010110110010101001; 
out28 = 128'b10010111101111101010110010011111101011110011111100000101000000010100100011010110001010111100001101110011101101110010000110010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out28[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out28, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100111101110000101101101000101111100101001000101010010101010011001010001000011000100111000111001010110011101110010011000101; 
out29 = 128'b01001001011000110110101110000110100010110000010101100110000000111001001011000111010001001111001100000010110000111100111100000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out29[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out29, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001101111000000101110101101110110001110011011010011111101101111000110001010100001110000011011100010100011000110101011000001100; 
out30 = 128'b00110101000110101000000000100111110000010010110101110101110000011111100110010011010010111001101001100110100111000101101010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out30[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out30, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101010101000110111010101110001100000101111100111011110001001100011001001010100010010000101111110100001010101101001100111111; 
out31 = 128'b00111011010101011101010010111110011001001010110011111001000000111101101010100100010101001101001110110010001111001100011010001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out31[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out31, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000011010110001110001010100111101111101011011001001011100010000100000011000001101010011010000000111010010111001111101011001; 
out32 = 128'b11000000100000101110000110000100101000010001000000001100101011000101101000111000001110010101000001110000010101000110110100101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out32[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out32, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000110101011111100011100110101101111010110011110001010111011000110111101101000001101111111001100000101001100100111101100000; 
out33 = 128'b11010011001111000111010111000011111111011110100111000101001011111100100001011000111101000111000100011010110010001011001100001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out33[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out33, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010010000100111011011100110010100100101100100101101000100000010110011001001100101001000011000101000011110101110010001110000; 
out34 = 128'b10010000010000011101001101111010001011111111111100010010111100011101101010100100000101101110011010010011000100010011001111110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out34[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out34, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110000101111111100100110110001011100011101010111001100101011100110101100100000111111000101101000100000101111111001110010111; 
out35 = 128'b01101011110001110100101111101001001101100001110011001000100011111100000011111000110001001011111001011110110011001001101101001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out35[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out35, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110100011100010000101100110000010101010010111111100110110111101010001011110110111000000110001000100110011111111001001110101; 
out36 = 128'b01001110000001111110111100011001011101000100010010111001010011110101111111111000010010011001101101111101111101000001101010111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out36[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out36, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111110010101010001011000001111100000001011111110100110110111011100111110101001110011001001011111110011101111000110011101010; 
out37 = 128'b10111111101011110111010011100001001010000101010110001101000111011101110110001110001110100110010010101010101011001001110010111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out37[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out37, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110000000010111110110000101010101010110001100111010100110101110010000111100111001011011100101010100001101000001111010000001; 
out38 = 128'b00010010111110011100101001001000011101111001011101010001000110001001101011000100010110011110100000110001110010010000101111101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out38[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out38, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110100001110000010010010010001111001100011100010111011110011000010010011110111010000100001101110111001111100100001100110000; 
out39 = 128'b10000011111110100110010111101110100101111000100001011101111000011011111000011010101100100110010011111001110110101000110100011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out39[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out39, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011011001111101010110110010111110010110011000100110101111110000100001010101001100100111001110100011010001111001001010001011; 
out40 = 128'b11100011011000011111110100010011001111000011010111010001101010010101000111110001101011111010111100000001001110001110101001010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out40[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out40, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010011111011010000110100010011000001111101111101011111011111000101101011001111111110101011000110111010010001000110111001011; 
out41 = 128'b01111010101110010001111001010111011101010001101110011011101111000000110011111011011110001000110001110000011010011111000110001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out41[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out41, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001111100011110101011111101101000010101110101100101010110111000000000100001111101001001010000111100010111001100000101101110; 
out42 = 128'b01000110110111001101100010110011100110100011101000000000000110011011001011111011011101101000000011100100010011010101110100111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out42[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out42, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111100110001101111110010001011001110011001001011010001000001101011000000000010000110000000101011100101111101010110110001001; 
out43 = 128'b00011001000101111110000001100100011100101100110000011101101010110101111011111001100011001110010100110100100010110000011001101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out43[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out43, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101100100110100000111010111001011001101100110011111100110101110110101010010110100001001001010101010101111001010111100001000; 
out44 = 128'b00101101001110101010000011011100110011100111011001100011001001010110000111111110010100100011011101101110000011110101000000011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out44[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out44, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000000111101111011101100101000000001101101111101010001111001000001101111110001001001001001010010010011110000011000101111010; 
out45 = 128'b01111110101011111011100000101010010001011100010000000010001100001111010000111010001010100000000000011010100001100000010110001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out45[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out45, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010101000010011000011010111000100111100111000001000100010100111101111011010011101000110110000011111000011010010111001010101; 
out46 = 128'b10111110111001001111100011111101110110110001100001011001110010111010011010001101000001110001111111011011110001101010010011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out46[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out46, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011000111000110110000010110010010101000000001001001111010101001011101001011000110101010010011011010101111010111101010000011; 
out47 = 128'b11110011000000100111010010101100001110111111010010010000011101010101100101000011010110110000000101011110111001101100100101111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out47[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out47, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001010001001000100011010110111000001100010000001011111100001000001011111001110110111101010011011011000111100010110011100100101; 
out48 = 128'b10001001110000101111100010100000101111101010000110011111110001101101001100110000011011101101001100111001101001001100110011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out48[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out48, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111001000110000010111101010001110001011101110100001111111110110001100010110001110111000010100111011000000010001000111100101111; 
out49 = 128'b10100011110111110000011000010011100000000000110000010101111111101100011101000000000001111010101100011001011111000000100111011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out49[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out49, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000001000010001101100111000100000011000000000100001111101101110001011001001010000000011101000111000011111111000000101011001; 
out50 = 128'b11001010011100101101110011011101100111000001100101100110011110011001111100001100100110101110111010111100100101001010100111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out50[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out50, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011001000110100101110100000010011100011100001000010001100100010110011110110000001000011001100011010100111010010111011000011101; 
out51 = 128'b01100000111100000111000001010011100001100010110111000000001010101001011010001111110110110111011010100010101001101000100011110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out51[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out51, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000100100000001110110010110111010010011001110101000001111101000110111101011011101010010011001010101011000011111100100000101; 
out52 = 128'b11000100011011101101011110110011101001100000011011001111010100111000111000000000111000110111001101110001100101100000110000011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out52[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out52, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101101100110100011100001001101000101010111111100001000000101110001110110110100011110010000100011101011101010111101000110010; 
out53 = 128'b00010101000010011001100011100111111011111101110101110101100110010000111100101111100001011101000111010110011111111001000011111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out53[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out53, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111011010101101101101110000000011010010010000100111010010010101101111001000010010101011110111011000010010101010010110101010; 
out54 = 128'b10010110001011110010010001000101011011000110000011010000001111110010100101100001011000010111101101110100100001011001011010010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out54[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out54, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111000101111010110101011111001011111101110100101001110011110100011010101100010000110110000111110010111011111110100001000010; 
out55 = 128'b10110000001110010101001000010010001001000011110111101110001111100101110000110000001011100001100000000111111110011101001001001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out55[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out55, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000110001100110101100100101010001100001011111111001011000010010001011010111100011001010111111011000001001010000010010000100; 
out56 = 128'b01111100001000110101101101100111001110100110100100111111110111010010011101000111010001010001011010011111100000011001101000001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out56[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out56, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011000110010010000100011110011011001100100100001111111111111011000100111000001111001111101111000010011110101001000110110111; 
out57 = 128'b11001100111010010000110111110110111110111011001010110111100110110101000111110001101000010110000111111001010110001100110000110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out57[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out57, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111110101110010000010111101111001001101001100100000011011111111110110011110100010011001010010100110110011110011111010100011; 
out58 = 128'b01010111101010001101001110101011000011000101011000011101110000000101011110110001000111101101110110001110001110001011100101100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out58[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out58, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000001001111011001011110111101100011101001011111100110101011001111010101110110011011000000111110111001000011101101010010001; 
out59 = 128'b11010001011011110100001111111000010100001101111000110011111111110100011111100110010111000000110110110000101101010101000111001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out59[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out59, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011111010011010000101101101110011010100010010100100010100110001010011100010011111101010110100110110000111101010101100010101; 
out60 = 128'b00010101011001000110011110001000101000100001101001110101011101100101001101100001110000011001011001011101001010111101111010111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out60[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out60, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111101001001101110011001101010001110110111000011010111011010001111101010111001111100111101001111010101101001010100111110100; 
out61 = 128'b00000100011001100011101111001000111001011100100101000111011101111010110110001001001110001101000000001000001001101100001000111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out61[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out61, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111101111111111011111001001111110001010111010100100010111101110101101110100111111011011010110111101011101110111011010110100; 
out62 = 128'b11100111000010111111010010010111011101010001111100111110001000101110000011001001000000001011011011000110100101011101010010100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out62[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out62, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100101111000101001010110010000001101011101101101010101000101100000101010011011001011111010011010000000000000001000000101111; 
out63 = 128'b11001101101000100010011000110001001111110110111100111101111011110010100010000001001010100010110011100010111111101111101000110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out63[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out63, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110110111001010111100011000010001101011011000100011101100010110101000010101011011000000110001100001101111001000010010110001; 
out64 = 128'b01001000011111000011100010010100101110101101001101101011011110111011111001010000100100100000000111000110010100001100100011011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out64[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out64, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000011100011101100111011000111101111110101010000110011110101010011101011001101010010100010110011111011101001110010111011011; 
out65 = 128'b10101100001011111100010110011000011111100000001111111111011011001101011001100000010001111110010000010111100100011000000111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out65[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out65, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001110111000010000110110010000101010011111010010010001001100111110110100010110010100011100101000110100101100010110110011000; 
out66 = 128'b00111001101101011001010110110100010101100011011110000011010100111110110100010111001111111101111110000110100010100101110011011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out66[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out66, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011000000110100000101011101101000000010111010110010111000001110011100110001010111011101010011100101100110100110010011100101; 
out67 = 128'b00110000100100001111011101001000010111001000000010111100110101010011101010101010001101100010011010101110111101111101010111110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out67[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out67, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011001111111010010010011110111101011101111110001010000101011111011101101110000100010011111100000010010100001010100101101010; 
out68 = 128'b00001100011011010011100101000000100110001101110001011001000001010010011001110000001000001111101101001000111100011111100110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out68[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out68, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010110111010110100000101101010111101001101110110111010011001001010100111000000011010010011010101110000011000111001110101010; 
out69 = 128'b00111101000101000011000000110101100010100110101111010011111111110100001110001000011001001110110000011111011111101111011000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out69[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out69, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100100101110010100010010100010011110101000010110101101010111111100000101101010101100111001110001011101100001111110011000011; 
out70 = 128'b10011001100100010110101100100100110111011100010010010010101110101000011100000000001110011111010111101111101001010111101100111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out70[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out70, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111110100010000111110010011011100001101001010111001010110010000101100000011010100101110100000111001110000011000000001111111; 
out71 = 128'b01111000010110011111101011011011001010000001101001111001010011011100010110110101111110111001010111100110101000100011010010001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out71[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out71, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111100000011110111000101011111101111010101011010100010001100011001010001001100011111011000111000001011110010011001000010010; 
out72 = 128'b11001110000111000110100101100111001101100101001011100111000100011110111010101000011010011101011100111000100000111001100100111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out72[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out72, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100011011100101010111111100111111100000010101000111110000011101110100100011101101101010100000001011000010110101001000000010101; 
out73 = 128'b00101110001110010000100000101110010000111101000001001100011101101100011100101000011111011001011001111101001011001011110001001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out73[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out73, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100100011001111101110010001101111000110101111101011011000010001101011011001001010000110000111100100100001111010110011000010; 
out74 = 128'b01100111010100001001110111111110101000101001101010001011110101000001110100001111100001100111000001000011010000100010101110011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out74[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out74, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001100010111110011100010000110110011001001100100010001001111010100110101010010010101000111000101011111011100001010000010001; 
out75 = 128'b10111101000110000100110001100000010011100111001111110101011010111111100000001100100101001001101101110001100110100011011101111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out75[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out75, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101001010111101101100100001101011100111100110100100001100000111111010111010100000011011111100110100101101110000101000000011; 
out76 = 128'b01100010101110100100010000000000110001100110011110111101111100100001011001001100101001000100110110001110110010010110010000011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out76[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out76, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001000010000101101001001110000110011100110110101110001110010100011000000010001010110110001101011000101001110011010111101010; 
out77 = 128'b00010100011111100101110110110101000001111011001000101010110001100100101001010001010011100111111111011101111101010001100111011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out77[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out77, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111110001011111011110000001001111011011000001111011100010111111111100100010010101100010111001011001100011101111000111011000; 
out78 = 128'b10010000001010000110001100001100101001000100010101111011010111010001111000101011110001011100011010110111001011001101011010100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out78[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out78, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111110100000010010010110000001010010001001101110101111100011000110101010100110001010001101001011111010011110001111011011000110; 
out79 = 128'b01110101101101000100001001111111010111110000100111111010010000000101100111011000001011001101111010010010000010111100011001111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out79[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out79, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011101110000100001101110100100011001000000010111111000010001101010110111011001110000011001001010110100001010001010000111010; 
out80 = 128'b11111000101111101111100110101110101011100101101000110101000111101110111010110011111011001100001110111011011011100000001011100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out80[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out80, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100111010110111010110111000100010111000101111110101111100110100100001110100101111100100110111100100000110100110111110001001; 
out81 = 128'b10100110111001110100111010010001100001110010001001110000011010000000001111100010111111001000010100010101000100111010111101100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out81[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out81, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001100101011100011000110101101001101001100110101110100111010110101011011101011110110100001011110111100010001000001000010111; 
out82 = 128'b01010100011001100111100010101101110000100101101100000011101110111010110110011111100111011100010010010111001010000010010011101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out82[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out82, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011110011000000010100011111000011001101001000011010010010110001111101110001110100000111101110111110010010011110101001001100; 
out83 = 128'b11101001000001011000010001011001111000010111011000011100100100101111111111111110001010110001101101100000010001100001010010100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out83[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out83, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010101101010100110110100110110011000100110100000101100000010101110111100001110001100101100111001000000011111010001110101101; 
out84 = 128'b00100000101011101010111001110101101000100001111001000101000100110111001101011010001011011001101110010110110000001010000100111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out84[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out84, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100000100011101000000001010001101011000110010101011000111100110001001110110110011001011010001101101111100001000000100001110; 
out85 = 128'b00111101100100101111101100100100100001111010110010000001110111001110010010001110111110101010001010100100101100001000000101111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out85[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out85, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111010110000010001100001010000101011111111110011101001110010000000111011001101010001101001110010000110010111111010110000110; 
out86 = 128'b10100000101000100101110111001000110011010001111011111101111011000110110011110010101111011001110000011110011001111001000101100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out86[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out86, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001011000010110010010110100111001000101100101101010000110001011100111100011010100111101000101100100001000100000101010011000; 
out87 = 128'b11001010110100110010011110101101100001000100110000111110101000000010101101001011001101110011111011111010011001010111001110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out87[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out87, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111100010010110101010101101011101111011001000010111100000011011101110110000010000000101100000001011100111010110011110111111; 
out88 = 128'b01111110101001010000001010010100101000100011001010011010111110011000001111001011010111111111100111101000001010010000111101110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out88[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out88, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110011000000111111000011110011100000110100010101011001111101110101011110111011110001110010110010001101010010001101100100011; 
out89 = 128'b11101111011010111100110001111101101000101011010000010011000100100101011000010011000010011001011011011011000111100110001110001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out89[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out89, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101010000100011001101010111001011111111101010110001100010101011001011010010111010110000000100010000001111011110100100000010; 
out90 = 128'b00100001110000001001111101000110011101011011010011101110011011111101100111010110111100011010011110010110011010101001001111010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out90[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out90, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101011011010001111011100011000111010011101111100111011000111011101000111000101000011001100001011000110100000100001000101110; 
out91 = 128'b10000111011000111001111011001101010001110010000010111100011100010011100101011111110000100110100101101000100110110101010011101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out91[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out91, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011001000111110010010111101100101001111100000110010001101001011010001111000011101011010010100011010011100001000011010001001; 
out92 = 128'b00011100001000100011000000001110000001000011011000111110110100110010010001110010001011100111101101110011011110001101101001010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out92[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out92, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001111111010110010011011000101101100111101011011100110100111101101110000111111100111110110110110000110110110000111000110011; 
out93 = 128'b10001001111010011000010100100000110110100111111110110100000010010100100001011001101101110010011100001100100111111101101001010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out93[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out93, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111111010011011001100000101011010011111111111001011111111110110011101011010110101111010000110111011111010111010011111100001; 
out94 = 128'b01010111111100001110101101101100101100101110011111000000001101101101000111010010110011011011111110001101000101100000110001000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out94[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out94, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010100100111011001101000111110001100110011010000111110111001000110010111100111000000011000011010011010101111001111110110010; 
out95 = 128'b01111010100000011100100101000110001011100110010100110001110100100010101010011101011100001111100101110110111001011101001011100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out95[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out95, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001110111100110010111000111110111001000010010111011110010111100100001100011110000111010101001111010110000110000101111010111; 
out96 = 128'b10000011100010010101000110111001111000100101011110010000011010010100011000110110001011001101011010000111110100111100000110110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out96[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out96, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010100111101011001110000111100011100010100100101010101011100100110001110100010001100111001101100011111101111110011110101100; 
out97 = 128'b00010110011011111110110011011110000010011000101000101011001111110110100110110111001110110000001010101111001110100100000110110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out97[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out97, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011100100101110011000011010110111000010011110101111111000001001111101110000100100110101000111010110011011110101001010111101; 
out98 = 128'b01110010011010101100110000100000101010110000110010000011111111011110100101100000000010011100001010111011100110000101110101001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out98[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out98, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001010101100001010000011101000010101010101001111110010111000101110011011000001000011101000101011111010100000110110111011100111; 
out99 = 128'b10000011001000101011110001110010111110100001110011010011010101000001110010001100111001001111101001001011110010010001100011110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out99[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out99, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001010000111100000100111100001000011101001000010100001010100100100010000111110100101011101100010110000111100000110110001001010; 
out100 = 128'b00110010100111111010111110011111101011111000111101111111110101111101100001001100111110011000100010000010010001000001110110110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out100[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out100, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010011111001110101110010100011100100010111010001011011111000000100101000010000110100101001101000011010101001101101010101101; 
out101 = 128'b10011001010010010011001101001011100001100100001111111001001001001100011111000100010011011101011110011011000111000110000111111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out101[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out101, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101111110001001001010001110100101011000011101000001000010100010111111110100011001100110000110111001000100000000100011010011; 
out102 = 128'b11110111011010110100011010001011010111001001110110111101111110011100100011111001101100001101001111111111001110110001111100111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out102[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out102, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101111000100010010011010001010001010111111101000010011010110100010111110010110001110100000101111011001100011110011011111110; 
out103 = 128'b01000011100001000011110000000001001110000101000010001111001001101011011111011000000100110100001101111001011110000100101001001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out103[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out103, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011110010001010111101111101011100111111111000010010011111001001001010010111011011010011011111001000110000101100010000010011; 
out104 = 128'b10110111011110010011000111110111111010111000010110011110001111100101011111010010010110101001000001011000100110111100101010110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out104[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out104, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111101001001100100000000000010000100110011001000010111010100000110101010000110100101111101101000000011111011000101000110111101; 
out105 = 128'b00011011001100000110110111000100110001101000010101110011100001010100001001100100011111001000001100001110101110111111010101111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out105[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out105, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001110111101100011010100000111001000000011100111110000001001110001010011100111110101110110110110011100110101101101111111000; 
out106 = 128'b01110111000011101110000000001000100000111101000000111010111101000010000001111111101100000110010100010100111110010100001000111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out106[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out106, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100111010111100101011101111111011010010111101110000111111010111111101010010111101101011011001001001000011011011000001111010; 
out107 = 128'b01110011100110110100011101010000000110101111000100110011111100111000100101000110000011011011011001100110001111000100011000011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out107[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out107, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000010010001110001100100100000011110101010011100110011101011110101000000000011111111010101101101101001111101110001110100001; 
out108 = 128'b10001010010110001101110000011111000110010000000011101010101111000001100101101011001110111111001001101101011010011010000001001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out108[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out108, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000111010111000001001010011010011111101101101001000111001110100111000111000101000110000011101110010010000010001001111011001011; 
out109 = 128'b00001100010100011100011001010011000000000100001011100011100001001010001101101011111110100000110001100110001010011111000111111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out109[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out109, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110101011011110001001010010111110110101001110000000100000100000111000001010110101100100010111101110010100100011010110011111; 
out110 = 128'b10101101000000000001011000001000011100011110100111000001011110011010001110110100111011010000111010111000111111010000001010011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out110[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out110, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000100000001010100110011110000110110100000100111011011111000011111010000010111001101100011011101110111110100100010010000010; 
out111 = 128'b00001101010100001110010110100111110000100000101000000110010101110001011010010111000100101101011110000110001100101011110110001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out111[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out111, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110000111111000011001000101110101111100010000011111100000000000100011111100000000100100000010001111101011010100001110100000; 
out112 = 128'b00010111100100101011011000111011000101100100000110101111101100000111011110111000001101000000110100111101000100100101100010000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out112[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out112, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011000010000010100000000111101000110111000011110010101000100101100010010101111000001110101100101101000010100010100011010001; 
out113 = 128'b01111001111101100001001010111010000111011101101011101010111100010111101000011010111011010111001010010111111100010100110001001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out113[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out113, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111111011000001101110100101110111001100101011100110101101000010101011010001101001101100001010110001110101101101011101111000; 
out114 = 128'b01000101000110000011111001111110111010100001110101111111111001111010111101101000101011000101010101100110110111000001010111001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out114[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out114, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111111011010110110110010011101101010110110001011010100011001010101001110011001011010100001101001000010101001011011011100000; 
out115 = 128'b00001010110010010101000100110011111101110000000010100111110011111100100000111001011000001011001010000000011101100001101001001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out115[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out115, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110010001011010010100010100010101001101000100110111111000101101000011000111000011011111010110100011011010100110110001010111; 
out116 = 128'b00100101011001110110111001001100100011111110000100101100000011100111101101011010100011100000111111111011110101010111101000001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out116[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out116, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111110011111011100100100101110001101010010010101110011110110011111010001100000010110101100100101111101001110000110011111011; 
out117 = 128'b01001100100010100111111000110100101011001011000011010111010011110011101101001100011101111101001000111101100001111011110110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out117[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out117, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010001110101111111111111100010011111001101100001110100011000110100010011101101000001110100110000111101111100101110111001101; 
out118 = 128'b01001011000111111101100111011100000010111010011001101010011111001001100111111101111111110011100000010101001111010111011011111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out118[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out118, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001001110110001000111110101000110100101110010111101011001001000101101001100001101111000101000000111001101000111001100100110; 
out119 = 128'b00110110010000000010100010001000111110111010000100001110111101001110000001000101110000101100010111111101010010111101101010111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out119[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out119, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100010000010000111000110100000001010101111100111101101111101011011101111101000100011000010101011011100001000111111101100011; 
out120 = 128'b10010001100001110101110101111001000110001001101110010110110011110000001100001111111011000111100111010010010011100011101001001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out120[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out120, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111010100110001010010111001110110001011010011001111000001110111011100000010111000000111101011010001111011011101001100100001; 
out121 = 128'b11110000101011100100110100110010100010000010011111100000110011111011110001000111001011100100110010011000001010100001010100000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out121[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out121, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011111101110010101001010000011110001100000101100011111100111110111001000101011100100100011111000001111001010011100011101010011; 
out122 = 128'b01010111101110111001011111100011000011100000001001011011100111111101100010100101011000001000100011110111001000010000010100010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out122[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out122, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011001110110101111111010110010111111101101001111010011110000101110101110001100001000101100001111101111001100100111010000110; 
out123 = 128'b01100000111010010111100100011100101110000101101000111011010111110110000110001101001111011010101100000101000111111111010100100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out123[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out123, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101000001001100100000001111010110000101100011011000101010101111101010100000011100010111001000100010001010010110111011111001; 
out124 = 128'b10001011100100111001110101010111101111111010101100100110010110010001110101001000100000100101101110010000000100111111011111111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out124[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out124, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001010000111011010010001100110001000101111100111010011001000100010101101111000100111010100011001110111111101000111100110100; 
out125 = 128'b00010111110010110000000110011011100101000011011011101101111110111100000110011100000001101001101101001011000011101111000011011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out125[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out125, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110100111000101010101000001011100101011001111100010110110010110100110110011110100111011101001001100110111011000100100110001; 
out126 = 128'b00001000100110100110000000111110000011100010000110110001011111011110100100010111001110001010000001001111110010100000010011111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out126[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out126, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011000011111010010010001110100101101010011110110011111011111010011010000001110010111111110111101101101011111000101100011111; 
out127 = 128'b01101100000011010101110010111111111011101111000110100101100110100000100110101100000000101100101100100111011110111111010000001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out127[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out127, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001011011101101110000110100100010011011101110011011111111011001001101111101011011001110100111010000100101100001100111001010; 
out128 = 128'b10101001010110010001011110111011000001100110111001011101001000010110100011010110000001100000111010110110100011100000010101001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out128[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out128, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111100011101000001101011001110100001100011110111110001010101111100011011000000100100111010001001100100000100001010101011001; 
out129 = 128'b10001110011111010110011001011010111101100001010001001010100111110010101110101011111110101101111011011101100001000011111001010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out129[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out129, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100011110111001110100110010101111001011101001101011110111100010000101000001100101101100101100010100010110000001100001010110; 
out130 = 128'b00000001011100111011011010111001001111110010001101001110110100001101000011000100000100111101011001010101011001000111001000111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out130[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out130, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100000000011110010101001110100110001110011010101100101101110110010010110101011011000100111001001010111011111101110011001110; 
out131 = 128'b00100100000000011110101000000001101111100110010100101101101110101010011111111101110101100000010111011111010100000001101101100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out131[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out131, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010101111001010111001111010110110001011011101010110111110111111010110100101001100101001010011011111111101111001111001101100; 
out132 = 128'b11001011101010010101011001101110011101101101101101111001110001000000011000110010101000001001011000101010001000000111001110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out132[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out132, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010000010011011001100001000011111010001011000110011110101010100100011001100001000010111100110000101100100111100101010101100; 
out133 = 128'b00101011001000111010001110100001010100010101011110010011011011101101111011111110011110010110010111001010111100011011111101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out133[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out133, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111010111000100111010000101000101001010101111101001000010010100000101111100101101010011101101000011010110001101111010100101; 
out134 = 128'b01101011101000110101000000110011001101011111011010011001101111000011101010011011100101010011010010111011100001010100010111000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out134[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out134, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100000010100011010100101001110001011001001001100101010101110110010000000011011101110100110110011101010101101100101111000010011; 
out135 = 128'b10001111011010001110101111000001010100000111000111100110100010010101110000000001000101001001101001101111111110010001111010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out135[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out135, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001100100011110001110001000000100111011110101010011110011101100011001001011000000001010000001100001010100101011010100111010; 
out136 = 128'b10000100000011110011101101100100111110001111010011111011011000100110110010000010111001111000000011110101000111101010100011111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out136[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out136, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111110011111011000100010000001000101111010110110100010101000001100101101111100001101111010111001000000000001111001100001010; 
out137 = 128'b00100011111110101011001110111100000100011100111110101010000000010100011011110110111100111011101100010110101110100000000111001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out137[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out137, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011010010100100110011110100000111100010100000000011001001001110010110001111011100101000010001011010010001111001001101101011; 
out138 = 128'b01011010100101110000101100110110010101111111100111101010111001000100110000101110010000010111111101100100010100110110010011001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out138[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out138, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010011001011010001000101010101111010110001100111011000101100100100100010101000101100100111111000111001011000010100100110001; 
out139 = 128'b01101010000111010101011011101101010111010101001000011100111000111100001110001101011010100001010100100111011111001011001110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out139[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out139, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001101101111110111000010011010001010111010110000100001111101101111101000101000000101001111111010000110110001010100010001111; 
out140 = 128'b11000000101010111111011101011001010010111110011110100110101010111111111111000010100010111111100101110111110111101110100100111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out140[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out140, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010110100111010100101010011110111011100100011101111011101010000110100000011111000000000000000100101110010011010100111101011; 
out141 = 128'b11100110101101111101111111000000000101001011001111101111001011011011100111110111011111100011101000110000111101011111010100100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out141[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out141, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101011001100001010010101100001111001000010001101010010001101111001111100101011111001100011111111111110001000110100100101110; 
out142 = 128'b01110110011111000100111001001111101011100100001111011011100110010011101100110110001101101110110111011001011101101100111001101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out142[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out142, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101110001001011100110111011010001101010010101000100001100000000100100010111111101010001101011101010010001110110101010011001; 
out143 = 128'b01000101001100101011101000100000100011111010111110000010101101100111011011011001101001101100111111100110000110001001001110100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out143[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out143, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010100011111011001000011100001001111001111101010110001000010110010110110011101000111110011001000110110010100100111110011011; 
out144 = 128'b00000101111011111000100011101110110100000111010110111100110101100000010000010110010001101001000011100001111100001100101110110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out144[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out144, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001001101001101111110110011001010011111101010000100101101110101000011000001010001001101010010110000101110110000001011100010010; 
out145 = 128'b00011110010110001101000110010111001010100000111111011000111001111111101100101110011010110101100110000110010000011001110001100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out145[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out145, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101110011111100101001011001011000000011100010110001101000111111101100011101011001000111111100110001111011101001101001010100; 
out146 = 128'b11100011100011011010000110101011111000111110001011111001010101010101001011010001100001110111100011010010011100001001100010100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out146[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out146, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110001001110000001010101011001101100000010110100111000011001010001011100100000000110110011010000011100010001100000010010010; 
out147 = 128'b01111100000111001011000001111101010000111110000110000001100100001111100101101110000101100110010100100101100010001000001100011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out147[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out147, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111000011011001100101100100111011000101011001010001100111000110000110001111111111001101110010010001001011010110100000000000111; 
out148 = 128'b11000111101110000110110001100011101101101101111010101101101010011011110001110111111110001011111011000000110011100011111101100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out148[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out148, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001010010011000110001000001001011101011010100011000111111011110011010110110010101011010110111110101000110010101011100110010; 
out149 = 128'b10100110000100011100000111000000011010110010000000011100011000010111111100110010110110100111011011100011111110011011000011111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out149[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out149, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010010110011110100000001011100111110010110000010000101100011011010110111111010011111101000111010001011001101101001010110100001; 
out150 = 128'b00001011100010110011001101011100011010100111100110010001011100000101010011100110000100011101001110101010010001111000000101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out150[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out150, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101011011101001100110010010100001111000011010101001111111100110111111111111110101100111100100110000000011001100101110100101; 
out151 = 128'b10111011010100100011010111100101001000101101111000010001110010001110110111011110010011111011001000000100001111011110110000011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out151[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out151, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101101001101011101111001011110000111110001011100011011011100100101111111011011010001000110111100101111110010010011101011101; 
out152 = 128'b00111101101010110100011010001110110001110001011011001011010010001111011011011010111010100111101100110000010101001111101110110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out152[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out152, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011111001011100111010100111111000101011111111001100110110110100100110111110000000010001110101011010010101111101110100100110111; 
out153 = 128'b10011011010110001111110001011111011010011101001110110100001101100000010001100100011101111111100100011001011010111101011111111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out153[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out153, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110111010100100111101000001111100010100000011110111101111110010101010111000101111000111100100010101001100011011100000001011; 
out154 = 128'b10100010111010010010100111000010110101110110001011011101110011101101010001100101010000111100100001001010101100001000100110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out154[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out154, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100000001100010100110100111100100011001100100100010000001011101011110011110010000111101101101101001001100000100000001000011; 
out155 = 128'b01000001111001010010010110011101011010101000000101111000001101101101111000011010001111001001010111010110000010011010110001011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out155[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out155, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100010001100001011001001100010111010011101011100101000111100101001010111110110001011111100010000111101100010110000001110000; 
out156 = 128'b11011101010110110101010101101001001110100100011110111011000110101100111110110000010110011001010000010001101111010100100001100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out156[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out156, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100011000001110001110110111110001101011010010111011010011011010101111011110101000100100000111100101111011101011011001000101; 
out157 = 128'b10101001111001111000001100001000000011011011110000011000111011101101101001011101000100001000001110010111110001000010111110100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out157[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out157, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000001100101111011010110110101001110100110110111010101011000101001101110011010100010001000010111000111011101010111111101111; 
out158 = 128'b01001010001111111011001011111101010010101100000110010000010111111111110111010101011000100101110001001110101011100001101101000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out158[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out158, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111110101100101000101100011100101111111110111101010001101100111000110000001110110110100110111111001010101110110111101111011; 
out159 = 128'b11101000011101011001110001111101000100001001000111010001010101001000000011110110001111100110010001100101000110010101010000110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out159[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out159, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100000000011111011001111001010101101100110101000111111111111100011001111001101101011101110001010000101101100001011101110111; 
out160 = 128'b10010010111011001011011000100100001000110010011111110100100010100000110110001111101101010100101100101111001101011001010101101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out160[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out160, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101001000000011010101010110000010101000111001010110000001011101101001011101110000101111110001110011110010001011010011000110; 
out161 = 128'b11101101001000000111001101111001100000111000011100011111011001001100111010010011001111101011000101011101001111001111100101101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out161[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out161, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011011001010000000101011001101000101100000010001010011010010001011110100101001010100100111000000010001101001110111011000100; 
out162 = 128'b10111101111111101100010010011111100010111001011011110110010001111000011011101011001110110011110110100110101000101001011110100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out162[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out162, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110011110110111101000100111111110110110010011011101010001100010111001110111110011101010111101111011011111000011110110111110; 
out163 = 128'b10010101001100000100101111100011011111101100001000111100011000110110000011000110011110110011110111010101010011110110101110010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out163[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out163, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010100101011001010100110011001101111001111010100001101000101000010011001000110101010110001010111000101101010011110101001111; 
out164 = 128'b01101000101111101110000101011001100011001001000011001101011111100000001100101011110101100100011100111111110011010001001100110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out164[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out164, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010110010111110000010001100111000101010100111101010001001010101101010100001100100101100101101101000110101000011100111000100; 
out165 = 128'b00111000101111010000101101010010111101001100111100100010000000110100111001111111001011111011100100111011001010001001100001010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out165[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out165, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100101001001011011111000001101011010101011110111001001011111101011011010011111110010010111110011001010000000100010010111101111; 
out166 = 128'b01000111101110111100001111000101001100110110000101111111111111101000111001110111100010110111110011001100010111110110110000000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out166[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out166, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110101001001110111001001011111010110001001011001100110011100100101101110010110101101111111001000101110011010011001100011000; 
out167 = 128'b11010000111111001111001101000011100110000100111010000000111011111001101100101100101011110111011111100011111100000100000101111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out167[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out167, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011111010100010001001110000101000011011101000000110011010001011101110111110101110001100000110101000100110111101101001101001100; 
out168 = 128'b11111100001000011110100111110101110011011001000000100101100100001100000000100010010011000011000111001010110000000100100000111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out168[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out168, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000000010101000110000001101101011111011111100010110101001001100001110101001010100001010010101000011111101010101100010010101; 
out169 = 128'b01110011101111100000110001001100010011110110111011011011010000111101100110011100111101010010110011000001111100001001011100100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out169[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out169, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001001011001110101101011010111011101111110011011111110111011010110001010110000111010001111010101001001000010000111101110000000; 
out170 = 128'b00001111111000110001000101110010001110000010110000100011011111101100101000001110111100011110110011001100111111000000001011110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out170[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out170, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001100000101001101110001011000010101011010110111000111101101110111011111100011110110110110100000011110011110100011001100001; 
out171 = 128'b01111011100101011101000111001001010110001011110000010100011011011100111001001101011001010100000111111101110001001010110101010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out171[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out171, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111111010000011100010011001111110111101010001010110111011111011000110100011100100000100010000011111110010110000001100111001; 
out172 = 128'b10011100101110000111000110011110001111100000111011000111011101001101101010110100000011101001100111110011001001110011000001010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out172[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out172, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111111101111110010100001010001111100110110001110101110110011001010101110000100001100011001010101001110111111101010010000100; 
out173 = 128'b01011101111100100000110100011001110010011001111010101011100101101000011000000100011000110110000101101110000100010111110100100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out173[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out173, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101100111110000101001010101110011011100001011111111110000011111010110000100100111110010100110110011000010110100111110010010; 
out174 = 128'b01111110010011111110011010010001000001000111011000100000100000110101110111101010111100100110111101001101011011100010000101000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out174[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out174, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101010110001110101110000101011111010011100000100111001110100110100011100110110000001111100111110110011011110111001001111100010; 
out175 = 128'b11001101011100111101001100110110000000100111000101100000000011011100011100100000001100111111101011110001000001011110101101010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out175[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out175, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111110100011110000111010010100000111101011100100101011000001110001111010011010010000001110001001100110010101111100100101111; 
out176 = 128'b00001011010001111100011101111101110011010011111000011000011101111000101111111000011100101000010000110100010111110010000110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out176[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out176, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011100010011000111100000100101111100101010001001001000010001101011001111100010110101101111100011100011011011001010000010101; 
out177 = 128'b01000000000011101110001001000001011000111111010111010101001010100101001110011110001011001110100010001111010100010111011110000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out177[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out177, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101011101000001110001000010100001000111001101011110111011111110101100010101111101100110100110010101110011111101010000010111; 
out178 = 128'b01000100010010001001111001111101010000100100101011101111101001100111001001000101111010110010011111110100100100010011011110101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out178[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out178, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010010100100110100100110110000100111000100101011011000010101001100001111110000011000010011000100100011101111010111101001000; 
out179 = 128'b10101001110010001011100110011100110000100011100001010000001110100001110011111100011000110001101111101100001101101101011101010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out179[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out179, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001101000000010101101101111000100111001101001111110000001011000101000101001010100111101100010100111001111011011101100010000; 
out180 = 128'b00000011100010001011001110001111000011001010001111110110010010111111101111000000111001000101101011001000010100100000010111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out180[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out180, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100010110010011010011011011100010000011001001111010010001011101111100011111010000100000110010101100001010100010011110011011; 
out181 = 128'b10011110001110111000111101010101111100111010110100101000111101111100100010110101110101000010010001111111110000110111100110101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out181[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out181, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110010011101000101011111101001011010001011110000010101011010000001111011110111001110111111100001001010110110111001101000110; 
out182 = 128'b00011001101111111101101000011100000111110001010000100100011110000010001011001010111101111100001001111001001110101111011101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out182[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out182, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110100111000100011000100001111000100011010011110000000111000101100110010100001000001111011101001000110011001111110101110001; 
out183 = 128'b01101101101010100111011001011000100001010001011100010101110101001110001100010010000000111100101100110101100100001100010101111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out183[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out183, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010000001100001010110000011000010011111000111001011010010110111000100000100001110001100000000011001100111101011001000001000; 
out184 = 128'b00010010111000000001010001110000111000110111000000000011010101100100000011111010101010000100110000000101001110001101010011101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out184[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out184, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001011100001001010111011100100101111111000100110100101000111100000111111100101001111101011000011110010000101001110011010000011; 
out185 = 128'b10111110100001010111100101000000110001010101111110011001111110010101010100110110101001011111011101100011000100110101100111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out185[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out185, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111100110111111001000111101101101000000100111100100110100001100110000000001011101000100111101001001101101101001100110010000; 
out186 = 128'b11101001101000110101111010011111000000011001111000011100011101100111100110011011000100101101110011101001100101010011001111101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out186[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out186, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011111010011010010111110110001100111000101111011001001111111110001010011110001101011110000110000110100010000000110001100011; 
out187 = 128'b00010110100011011110001110010011001111000111111101001000101111100011000111011011011100101110010000101101000011101001100110110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out187[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out187, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101101100110011000101010010001001010001001011001000110010110101100100011111110010110100100011100001101010101001010101010110; 
out188 = 128'b11011010100101001011101000011010010110010100100001010110010001001000101011111110001011101101010001011101010101000110010010001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out188[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out188, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100000100111110100100011010100111010110100101100110111110000010000110101010101100100001000101111101101100011010100101110101; 
out189 = 128'b11110010110110110101010110110111111010000111111011110100111011011001100101100011000000111010100000001111001100011001100010111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out189[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out189, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110110111111000101111110111110101011100101101111010101111100000100011111110000111001101110000110100110110111101011110011000; 
out190 = 128'b11110111100000000100110011011111011101011010100001000101110101101001011000110111110110000011000111011010000000111001101111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out190[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out190, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010010110000101101000111110101101100101001101010010111100010101011010010011001001111110100111110010110001110010100101001101; 
out191 = 128'b11001011010100110110100000000111111011011000010111011000000101001111001110011000111010110010101011000001111100100110110010001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out191[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out191, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101110001111001000101010101100101100100011111100100010011000111001010000011011001000000110011010000100000110011100001001100; 
out192 = 128'b01001011111101111001001100000111110011001010000010001010010100001101110101110001101010001100010011011001111011011110100000001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out192[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out192, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001010101011011010100110001001111001001001110111011111111011111000110010011100010110011100010101001000000001110100111001011; 
out193 = 128'b00000011000101011111000011100111111000011110111000110010000101000101001000010010100010101001111111001000111111001110100101010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out193[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out193, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000010101110001111001110111100100101001110111011111010111000001001010011000010111000000010101110100101011011010000111000111; 
out194 = 128'b11101111011001101111100111000000001011011100111001110110001110100111000010010110100010010100001010001001111000100011000010101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out194[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out194, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111100100000111111010111100011000101110111100010101111111001010011100101011010001100000100001000101110100110100101000111110; 
out195 = 128'b11000100000110100100101011101010101111100101000101100100010100100110110110011000111011101000011111011011101111010010110101000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out195[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out195, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101001101000100011111111111100111011010100111011111110111001100101101110101111111101000111111010101000100110001001000011000; 
out196 = 128'b10111000001000000110000000101111001100101110100101100111011010100101010001000000101110111000110110011000011101110101100001000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out196[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out196, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100011011111001101000100010000001000111000010011100011101010000001001010101101011010111001001001110111100111110001111011100; 
out197 = 128'b10100110100111001000011000101101001011000001100001111111110010010101011111010111011101100011000111011110101100010100100001010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out197[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out197, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110011111000010000101000110100000101011000100100011001111101111010001001010111000110111001010000100001010110010110001011001; 
out198 = 128'b11011010111101010010010111010101010010010000101000100110110010100000001011010000000001011100111010011100100010000010101101001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out198[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out198, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101101010100111011101000000010010010100101010000000100101100000111011011001110110011001101010111000011000101010111011001011; 
out199 = 128'b10011001101111000011000000101011111110101011100101100011011100101001000110011101000110001100111010001010011011011110000111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out199[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out199, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111001001111000001000010011111110101110000000000110101101100110110111111001011000011101111110011110111000100001000110011111; 
out200 = 128'b00100010111010011101000000111001100100110110010101000000011011110011111001010001100110111011101101111110101100010101011100111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out200[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out200, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101101110010110000111001000001011100010010110011011101010110110001101011000000011110111100110010110101000100011010010111001001; 
out201 = 128'b00101111110000110111111101111010010001000010011010111100010010000111011000101000010101010101011000111000010101011001000111101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out201[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out201, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000100011000001011101100000001001011010001100000101000000010000000100111101010110010010100110000001000101000010010100010100; 
out202 = 128'b11011000110011010100110101001101110111111101011100110000101001111010100010100011010000000110111100110111011110000001100100010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out202[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out202, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000010010000110101011111110111100101110010010111101100011001110011010000100010111001000001111010110101100011011001100011101100; 
out203 = 128'b10100101011010110110001101010001011111110000110001010010101110101001101111100101111101011110000001111010101100110101100011001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out203[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out203, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000101000111110100101011111110101000010000010000011011100000101101011100001110011111111111100100001010111001110001100001000; 
out204 = 128'b11010100010000100110110001001011010110000111001011000011100100100001000111001111011001001100100011101010000001001010001000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out204[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out204, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010001111111110101100101011011100100001001110010100110011111111110111111011000100111110010100000100001000110100011010010000; 
out205 = 128'b10111100101011110011100000011001110001101010100011011010111011001000001010111001111100011111010011110011010000001010110010111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out205[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out205, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000000100101011111001111011101001111011111000100101101010101101000111101110111110100101010101000011100001101000100000110101110; 
out206 = 128'b01011000011011110100110011001111001000011101010011111001110010111010110100110111100111110100011000111100000110010100110000111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out206[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out206, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110010111110010001110100011111010010000111111000110111011100101001001100010011000110111011110111101111011101110111100110001; 
out207 = 128'b10111111011100010110000101100001010011100100111111010001011011100000110101010000100011100111001101110110001001110010100000001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out207[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out207, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110010100000110100010001101110000111011111000011111101010111110011011000111100111111111110101010110111011100001100011111101; 
out208 = 128'b00010011000111101011101001010111011000010100011111010100100001001111110111101011011000011110000101001010110110100001110011110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out208[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out208, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101001111001110011110111011011000000110101110111110000100100001011000001000010110001100100101100101110111000010101010001101; 
out209 = 128'b01000110011101010101110110111000111110000100111011100111110010000110100011001100000101110101010010001100001001110001101011001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out209[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out209, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001100100011111001000001001010001100100000100101110000011000100001001000001000011011101110111000011000011010100100011111000; 
out210 = 128'b11000100111001011111001010110001110000010011100001011100010110010010010001000101101111000101111110101110000001011000010011000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out210[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out210, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011010010010100000101111101000111111110110000101010001010100001101110111001101101000111100001001010110010111100110011100110; 
out211 = 128'b01100100000110101101111110011010000100100110100111111110001001001110001011100010110011110010110100111110111100100001011100000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out211[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out211, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001011010101110110110011000010111111100001001000011000011011001001111100111010010011110101000100011101010110010001100000001100; 
out212 = 128'b01011011011000101010110010100001000001100101100011110001111011101000100011110010001000010110111101110000011001101111111101100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out212[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out212, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011011101100110001100100000100010000010100101010000111100001110011000101101111100110100001111111111001010011000111001011011; 
out213 = 128'b01101110100101111100100010111011101010011111011110111011011111100000111010101101010001101010001100111000111001000111001000010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out213[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out213, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010101011100001110100011111001110001100101001010001100111101010101101100110010011101111100100001100111000111110111111000110; 
out214 = 128'b01010000001011111010111110001100011100100110011111100010101010111010001111011001011110010011100110111001000111100011000001010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out214[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out214, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000100011101111010001001011010000110000010100000111011011110001001000011010111001111011001011001111100100010101011000010010; 
out215 = 128'b00011001100011101110111101011101110111010010000110000001010010000011000110011000001010001111101110001011001001110000000010010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out215[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out215, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111110110100110100011100011001111011101010001011111011010011111000010010101001101000100010110000110111101011110001011011111; 
out216 = 128'b00011010010110001101100011000111001010110000101100000111111101010100100010011010010110010100110001101111010001100010001110100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out216[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out216, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001000101000111101111001101111001000010000110001001100010110110110110000011111001100010010010101111011100110100100111100110; 
out217 = 128'b01110001111111001110111001010111010100001000010000010110011010010001110011100101010110101111010011011001111111100010111110111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out217[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out217, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000011111000110101101100011100010110010111111010111011000001010101110000111011000001110000000001010000111110011111100110111; 
out218 = 128'b11000100010001111010011001100110100000001101001100001100101010011110001101100111011111111100000110101101110001000111010111110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out218[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out218, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100010001110111100010111001110010011110111010101001101000110000101111001011100001000111100110101111101000100000000000111010; 
out219 = 128'b01110101111110101110100111010111001010101011111111110011010001100011101000101010111111000101111101011011011100001110111011111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out219[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out219, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011100111111100100000101000010100100111111101100011100000110110010001001010110100001010000010111100010010000100111100000000; 
out220 = 128'b11000110010101011001101110011000111110111100101110000001101011010000110010011110000101100000111000110100010001101111001011111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out220[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out220, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000100010110011000110010000011101011110000001100011010001111111011111000010011001110001000101000000100100110001001001011111; 
out221 = 128'b01101111110001100111100110010001001101001100011010110001100101001010111110011110000100111000101110010101011111000101110011000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out221[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out221, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001001001000100000101100011110000101101010011000001000011100011100100101000101110010000000001001101001100101001101101010011; 
out222 = 128'b11111100011111101010011111100100011001100111000001111010111001100010000101010000101011110110011011110111111010001011111001000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out222[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out222, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110011111100010101111101101101011001100110011011001111001100110011111101010010001110110111100100011100111000000110010111011; 
out223 = 128'b11001111011001101110111110000110101111001010000011010001110110010001110100110010001001011010100001101001010101111100110010010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out223[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out223, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101011010011111011100000010110010110010101011011111000111110101001100000000000000010111111100110110010100010001101111110100100; 
out224 = 128'b10101011110101010100100000000011010110000111000101110011100100101000001011100001011000010000111010000011000001011001011101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out224[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out224, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000011010010101111011001000011101011110100011111111000010011110100011101111100001001001011110010001101111100001101011001111; 
out225 = 128'b00000100010101010111011011101111100110100011010111000111111111110011001010101011100110111101011000011000101110101100110000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out225[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out225, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010111100101101100011000000011011000111100011010101001011111011011010011010110111110100001000001101000101110011110101101110; 
out226 = 128'b11001110000111100100101101000010101011100101110011011100010110110101111111100110111011011000101100011001100010010100100101000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out226[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out226, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010110110011011001111111100111010000110110011101010011000100111001110100101000000111111110100111001111110010111101111110110; 
out227 = 128'b10001101111010111111110000010100000000001111001110111011011000110001101000100011000100000100100001111010110001000010100111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out227[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out227, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001000110011000001010110010011011011100110011010110111000011000101001111011101101001110111100000101001101110011001000011101; 
out228 = 128'b10100010110110010000011111001000010010100000100101101111001111000101101111110010011011111000011001110010011100001000111111001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out228[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out228, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100101010011101100001111010011000001000010001100111100001111111101000010011011011100010000010010110100001001001101101001100000; 
out229 = 128'b11110111000110110011000100101111000100010101101011001010100011011101100101000011100111011110100111101100101111101110101001111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out229[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out229, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001111111100011010000111010101010111001001110111101010110110000100101110001100110001100111101011001000101000010001011010100; 
out230 = 128'b01000001001001011100101010000101010011101011000010110010011010000111100011100110101110000101011011001110011010100011001111100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out230[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out230, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101011101011100100000100000111000101000100010010101111110010110100001001000000001010001000101111011011111100101011001100110; 
out231 = 128'b00010100011110011000100011000110100101010111110011101110110110011101100111011110001010011110101010011001000000110100011000001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out231[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out231, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101000000010110010101000110101111100100110111101011010100100001111100001010000110110000001100111001001110100011110000010110; 
out232 = 128'b11110010001011111100101011011010100100001101010100011001010100000011011111010100110100100100110110011101111110110101110110011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out232[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out232, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001010010001100100010011001001000001011000001101001110111011101011101010101010011000101110101100100110110011101001011011000011; 
out233 = 128'b00101111111001010111000001000011011100100100011011111001111111000000011111000101101000110110110101111101111000001110001110000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out233[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out233, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110000011101111100000101001011011100010110000000001110000101010111011110011010110011011101100000001100100100010011111010111; 
out234 = 128'b10000010100000111101010100100110111010111110001010100111010000111100111001110011101100001011011100010110111110100010000010101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out234[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out234, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111001000101101011000011011000110010101000001100101011101101000000001100101100110000011010101010100110000100001110000101011011; 
out235 = 128'b11111000010010001000011010011000111010001111001110110110111111101000100011100100111010111101100110001110000110101001000011101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out235[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out235, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001001010011011011100101000100101011101000101111100110011001011100011010011100010101010011101110100000101100010101000010110; 
out236 = 128'b11100110010011011110011111100111111110110111110001101100000010000101101100110101010000101001001111110110101110100001001110011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out236[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out236, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110011000011011111100000100001011110000011010010100000000110000111110000100111100011001100111001000101110111000010110010100; 
out237 = 128'b10101011101010010100101011111101100011110000100011111000011000000001111011010110100111010100011111001010100000100111000010010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out237[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out237, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000011010010010111101111000000100001010011110110000110010010100100010000101011010101111010001001101001110011000010101110110; 
out238 = 128'b01110100110001011001110001011000011000111010011011010011100110011010101001000001100111111010111111101110111101011010000111110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out238[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out238, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000110010111000101001010110000011111100110101001111111001011000010111110100011111001110001001001011100111000010010110100010; 
out239 = 128'b01100101010101011100101001111010010011000000111000100000111101111001100111011101000000110101100101001000000111000010000001011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out239[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out239, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001010100000101110011001100111001011110100010111100100001011010010001001000010101000010010110110101010010011111001000011010; 
out240 = 128'b11101101110101101100111011110101101111101110011010011010011100110101010010011000011110010110001011111100110111100011010110100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out240[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out240, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111010110000011010111001010011001010000011010000111111011110100110010111010111000000100000000101111000000111010011010000111; 
out241 = 128'b00110111110111001111010101111100101100100010110001110101111010011010101010011101101001001100100011001100100010010010011010101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out241[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out241, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111101100011101000000100110100110001010100000001000010000101111001010011100010001000110010011000110111110010101000011110010; 
out242 = 128'b01010001001110010111011010001101010000011000101001101101010001110101011011001111010010011010011000101010001001111011000100100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out242[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out242, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101010000111101100111111011011101001111110001111010101111111111001011100100000010011011000010101001011101111011101111111101; 
out243 = 128'b01111010111111110000011101011011110101100011100100101010110000111000100011011000110110001001000101111010010110000101110000100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out243[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out243, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001111011000000000001001100110101001111111000111111111011101000110001001110011001000000101000110111110011010001010001111001; 
out244 = 128'b11100000111010010000011001101001101100101100000001010111100100101111000101111010010011111100000010101010011111111011100111001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out244[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out244, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111011000000011001110011000001101001101101101110110100110100100010001010000011001110101100110010101011010111101010010101010; 
out245 = 128'b10111111100011001110010110101001001000111001110101100010101100000111011100001001100001110100000000001110111001000101110000100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out245[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out245, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001100101110010011110111011100101001110000010111100110011100001011001000101001100100110100101110100011100000011000100000101; 
out246 = 128'b11011010100001000110101110010000111000101011101001001010100100110100001001110100011001010110001010001110010110111101101010000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out246[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out246, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000111001000001010010100010100011100011000011101011101100100111000000101001110110011010101010011010101110100110000010010001000; 
out247 = 128'b00011001000000111101100011110011011111001110110000001101110101111101110100011111111110101010010011111001110101000110000101011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out247[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out247, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100001101011010110010000100111110110010000000110111001001010110000111100101100100010101100110111101010101001010011100101000; 
out248 = 128'b10011110100101001111001110000110000110000101001111000111010010110010101011000110011010011011111000011000101110100011011101000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out248[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out248, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000110100010111111110111101111010001000001110111001000101111010001111100010010100000111110000110000110110110001001000001101; 
out249 = 128'b11011101000111110011110010001001110111001011011011000111001001111100111110010000101110100010000000111100100110000101110111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out249[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out249, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101110101111100100110101010100100111110010110111011101010101001100111001000010001111101111001011111001101110001000110100100; 
out250 = 128'b11010100101100101101011011001101000110000001101011110100100000100000000100000111111000111011111000101110010010111100101101001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out250[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out250, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000111110111101110111011101111111001100101111011111101011100111011111100100001110110101110000110000000001010010000010111100; 
out251 = 128'b00010111000111001010010100110101101001010111101111100111001111100100111110001110011011101010001010101011001011101100111101110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out251[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out251, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010000011101111001100110101010110010110000011011011101101100110011110000000111101011101001010010001010111011011101011010110; 
out252 = 128'b11010011101010111010001011000111100001110111110100101010000111100011110010010000011110000101011101101000011011000110001100110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out252[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out252, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000010101010000011100010001000000000110110000100111110101001000110001101100110110001000111001010100110111000101001101011101; 
out253 = 128'b10111100110010001100001001100100000010001001100001110110110100010010110010001101000010011001001100111000110101011101011110101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out253[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out253, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010000000001100001101000111000001101100000011100001000110010001100011000100110001101110001111011000011010111100001010010000; 
out254 = 128'b00010111110100111111110001110000011111111001111001111000010010011111110001100001000001010000010010010010001000101001010100100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out254[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out254, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010010111001000000011110100100101101101001011101111011000001101011010111011110110110000100001101000101111110001011101001011; 
out255 = 128'b11011100110000001010011100100010100110100001101111000111011111000111000011100100001110001001110100100000110011111101101010001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out255[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out255, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011000011011010111011110100100000000111011101101000101010001001011010000001101101001010011100100001001001100011001101001111; 
out256 = 128'b11011001101110011010011100010100011101101110001100101100101100000101111001110111111010101001010101100001100101011100100011111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out256[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out256, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110111010000000111001101110001011001001101001010001110011100100111100001110010010101011110000111010001011100000010111110011; 
out257 = 128'b00101110010100101100101000110100111000011100110101000100111100000101110010001010011111101001101000100101111111101010110000101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out257[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out257, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110101111100011000111110010110001010100100101011000111010111000110111111011010101001100101001000110111111101001100100000000; 
out258 = 128'b00001010011100101011001101000101000110110010011010011100000011101000010000010101000010001100011000100110101111111101010010001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out258[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out258, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110000100011100100111111010001101001010111101011110101110111101101111111111010010011110001111001110011110001000111000111010010; 
out259 = 128'b00111010001110110010111101000101101000100101011110000001010111110010010010011111000000111100000011011001011000010010101101100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out259[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out259, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100101100001000101100011010101011100110000011101001101110110111110111100010011101011110111111111101110111000111110010100011; 
out260 = 128'b00010111000001001001110101110000010100100101011111011000110001001101111101011100010100101101000001000101000111010101100001110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out260[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out260, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000000010101100000100110110110100001010110110101110111011000110010100000110000110100001110101100110101001101011010111110111101; 
out261 = 128'b01001010011010001011011000011111001101100110111101110101011010101001000111000010011011001000011000001110101000010110011110100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out261[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out261, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111101000101000000101001000000100111011000101011111011100100101001111101110110000101101111100001110100000101001001001011010; 
out262 = 128'b01110011111011100110111110000000011001110000110010000010001001101001111101111100101100111011010001001100000111110111010110110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out262[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out262, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010110111000010011110100110110100010100000111010110101101001011100100011010111000111001100110110100001011000010011000011001; 
out263 = 128'b10111010010110001000000010011111011111111100110100110011111101011001100100110100101110100101111100110101110111110001100000101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out263[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out263, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100110001100101000000100111101000111001010100011010111111101111101101010110000110100000111001111001110011110100100010101000; 
out264 = 128'b00110111001011001101001111000111100101011111011010000101111001001110111011011011001011110111101000010101111111110001000011011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out264[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out264, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110000101001110110110010100000001011111100101011110110011101011000110100101111000100001010110000101001100110100000011111110; 
out265 = 128'b01011010110101011011110000000011001011000011110000010010101111110000111000101111001001101010110011100011011111010100001011111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out265[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out265, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011110010001010000110110100010110011001010001010001100111111011101100011111001001010010010011000000101000011011111100001011; 
out266 = 128'b00010000111110101010100110001110110110100111011111111110100101100100111100100110101101111111001000000110101111010101011111111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out266[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out266, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001100011100000111111110110001000100001111001001011100000000000100011110001100010101101101001001010011111011000101110110111; 
out267 = 128'b01010001001100011100110100011001011010000000010011000101110011001101100010110010010111000001111110011001110000000010000111001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out267[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out267, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111001100101111111010111101000101011010011110101010011010010000101000000001111011110000001010011011000001010101001001111100; 
out268 = 128'b00001111001111001011001111011110011100101001010110111000001101101011000111000101011011101010100101001110001101100101011011100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out268[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out268, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111100001101001011100000101011000011010011001100110101100010000111100111001011110010111101000001001100011101011000000001101; 
out269 = 128'b01001101011100110011100100010101000011001111010100000010101111110110110000001001101001100001100110001110011111011100011101101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out269[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out269, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111011111011111001010010101000101001101111101100010001110010001100001000001100100010100001010101011110001111101010010001000; 
out270 = 128'b11000110110101010101011101011000010001001101001000011010110010011001001101000001000100010101110100000101001111010111101110101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out270[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out270, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000100001001010110101101000111010000110011010110111111010111101000001110100101111011110010100101100100100100011100100011001; 
out271 = 128'b00100001001011010110110110111100110001001110010100110100110100010011010110111011011010010000001011101010101101000011101100110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out271[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out271, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010111010011001011001101001010011010010011001011100010101010000100001000001100010011111010000000001101110000110110110110111; 
out272 = 128'b10110011000000111000011111100000100010000000000000010110111000001111011001001001001000110100101111011111110101001010111011000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out272[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out272, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000001010011010100110111000111001000001110011111100011100110010001101111100000100010100011000100001111001001101110111111010; 
out273 = 128'b00110000110101110100000111001100001000000110010111100010110101000000001100100010011110001110110100111110100101111001011111100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out273[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out273, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011010010101001011100100101111001110110011010101101011111011010101101011011101110110011101111000100110000100111001010000000; 
out274 = 128'b11001010111011011110011101010010011010100100101101111001010110000011001111100011011101011011110101010110100110100101011010100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out274[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out274, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101001111100010000000011111101010101010111111011110001010110010110100101101111010110011101111000010100010111011010100001110; 
out275 = 128'b01110010011111010101110101000011011111111100001010000100001111000101100001000100101101101101010100001001110101001100110010101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out275[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out275, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000001010000000100101101111110111110000101010000110101001010010101110001100011010100000111100000111100010010010101111010000; 
out276 = 128'b11101001101101110000010011011100100111110010111111110001101101000010001111010111100000110101111011000110101111001101000011110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out276[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out276, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001111001010101110010011111111011111001100001101001110100100101011100111100101001000111010010110000010100101110111001000100; 
out277 = 128'b10011001111111110110011110001111111110010001010101110110101001110011101100011101011000100010101100110010010100111000001011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out277[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out277, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111001000100111101001110101010101111011100111101010001100000010101010010011110101100110110011000110000011101111000001011110; 
out278 = 128'b01101101110100001001111111110000000100111110010101000101000010111111101001011110010111110110111001100010110110101011111110100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out278[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out278, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011111010011100000011110010110010001010101010010100011000001011101111001010100100110001010111110101110001111110011110101101; 
out279 = 128'b11110110100101000100001100111010101100011000101010011010011010010111101101001001000111001011001010111001111001001001001011001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out279[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out279, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000001101000010110111101001110100001011010011000111000111100001101001110100110001010100011101000110010001100011101011011010; 
out280 = 128'b01110001000001000011110011000110101001100101111001001001001000010000111111010010111101001000100010111010001000100000100111010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out280[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out280, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000000000010011111100110100100010101100000101110101011100111000100011111011101011010011011000011011000110010110001111110101; 
out281 = 128'b01101101001010111101100100000011011100101100110010001001011101101011110011101111011101000010111111000111010111110000001001100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out281[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out281, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100010001110110010101110110001001111111101011000101100011101011110011010101111110011000100111001011010111011110000100001001; 
out282 = 128'b10100101000010111001001000100101111101100100001001110010000100010010110110101101001100111100110010010101000100100011000111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out282[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out282, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011001001110100101001011101001101101111111010010110101111110100111101110100001100100111011010000010011000100111100100110110; 
out283 = 128'b01101100110101011001011001001010001110111100100001000100110110100000001000111110000100011101000100000010001100011111101100000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out283[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out283, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110011110110011100011011001110111010110001001111100101111000010100110010101111110100001011111101111111111100111101001010001101; 
out284 = 128'b10101110011100100101101010001100111001100010000100101101100000011001100001011011101100001010001101010111100100100101111110101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out284[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out284, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001100110000010000101010011101110001110111000111110101111010100101100011110010111101011010110001111100100101001110001011100; 
out285 = 128'b00001111110100010110011100011111110111010000001100111101010111001000100010110111000010010010000110010011011010111100001100100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out285[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out285, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111101100101011101010001010011111110001110000110111011110111001001000111000000010000110011000100011000111000011111011000001; 
out286 = 128'b01001111100000000010011001010101011101000010100001000011111100010101111101010001111111111010110111101111110001010101010000111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out286[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out286, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101011000111110100001100101101001101100100011010011010001100110011110111111001001010101110000010110001101101101100111011111; 
out287 = 128'b10001011000100100001000011101110101010110010111010001100011000100111110100111011101010000010110011011110000110010011011111011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out287[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out287, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110001000100110000000101111110000000111011110100010001000011110001101000010000010010001111101100110000101010100001100101010; 
out288 = 128'b11001100000101001100101001000110111000010100001010011101000010011011001110111001010111101111111011110100101010010000010001011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out288[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out288, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100101110010110001001100010101011100101101000101100000011011110100000100110001001101110000110101011010011100111100010000111; 
out289 = 128'b01011001100110111101000011101100011001011011000001011110111100011110001000010011001011011100111100011010010110010110101011111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out289[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out289, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011011110110001011001111101110001111100101011001111011110011100011110010011000100101100001011111011000110110001110101010101; 
out290 = 128'b01011101000110000101010000000111000000101110011110110100100010110101010000000100001000000111011001111110111110111111001101001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out290[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out290, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110111111011100001001110001111110011101010011010001000110100010111111101010111001110001111000001110110110110100110111101000; 
out291 = 128'b11011101010101011101110011010011001011101011101010010000001111101011100110010010100100000000010001111001000010111011001101001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out291[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out291, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111000100010111100100010010111010111110101110000101111110011100110000110000011001010110101001110110101101001001100100000000; 
out292 = 128'b00011011001100001011011010000111000111011110000101110011011111010011011100000100010001111011101111010001101110011110111000110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out292[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out292, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010111001001100010100100101100101100010110011011110101111010111101110000100000100001001001110000001000101101011101010000101; 
out293 = 128'b00100101101010101010010001011110110010100101111000001101010011010110110011101110101011001011001111111111010100011011001011010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out293[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out293, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100101101010111111011111100001101100100111010111010010000101110101111110010100110000101011110001011010010011011110101110001; 
out294 = 128'b01010110100101101111001000010010011100000001010100110101100100101001010010001010111011011100111111101011011100101100011000001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out294[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out294, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001101000011110110111100011111000000000011000010101010001000010100100111000100101010010001001000110100001011100001010000001; 
out295 = 128'b00001101111100011000100011011010110101101100100001011111101111001000010111011110100101000111101110000111010110110101101111100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out295[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out295, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001110011111100110100010110000111101111110100110011111000100100100011010111110101011000101001101001101001100111100110111111; 
out296 = 128'b01111011001001111011110011100101001011000011011100110011100110101011110010001100010111011100101011111010101010011101111111110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out296[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out296, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100011000100100110101100111101100111000001000110110000110010010100011010100000011110001001001100010110110100101100101000111; 
out297 = 128'b11110001111111010111101101000010010100010011110100101000011010010110100100110000110101001101000011101100110100011101101101111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out297[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out297, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001100111101010110100101001101001111101101001001001100111001100011000001100010000101101111000011000110010001111011100100110100; 
out298 = 128'b01111111110010100111110101100000011011011001110100111010011001001011010100010001010101001100011011111101001011011000100001010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out298[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out298, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001010100000101010000011010100011110100101010101101011110000011101100010011011010010101001010000110011001101010000011110111; 
out299 = 128'b01000001100010011011100101000111110111001001000101101111100101000100001100111001000110111111011010110011000110101011011110101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out299[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out299, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010010101001000011100001001101000110110110010000001100110111010101111111001011100100010101110110011101101010011001000100000; 
out300 = 128'b10011111110100101100000110011110011101011100100001010001011110010000100011101010110000111100101010000111001101110111000010001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out300[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out300, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010011010001110110110100011101100100011011001111111001001100101101011100010011111000111010010010100101011100010111110010101; 
out301 = 128'b10101111110110111011101100000000010111010100001000001100000111001010110011000011010000101000101111011100010011100111100111100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out301[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out301, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001101000110110111110111000111011001111000011110010110001011001110011100000000010111100110101011011100001000100000111000110; 
out302 = 128'b01101010110101001101101000010001101101011010101001001111001000111111010110110110110111000101101101001111100000100011000001001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out302[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out302, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100001000100110011100010010100100111010111001111010101111101011101000010100011111000100111000010001110010110101111101110111; 
out303 = 128'b00101000001100111000101110110011110100010110111001101001011110000100100100111001010001001100101001011010000000000100101011101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out303[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out303, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111110100001001111111100010011101111001000001001110101110010100010101001010111010010000001110001100111101010110101110111110; 
out304 = 128'b01000101110010000000100001110000101100010111001101101000001100100111010100011101000010110101010100011100010001101100101000001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out304[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out304, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101110111001000110110110111101010100100000100101101001000111001001110001001010111101001011001111001100110010010101101110100; 
out305 = 128'b10100101110010011100111010010000100100001111011001000000000111001001111110011010001011111000000010000110000110010110100100000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out305[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out305, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001010111110101001100111011010001101001011010100010000111001100010010001001000111100010000110101010001100000000100111101101; 
out306 = 128'b00011010111010011011110000101100101111110100001101010101001011000110110111111101111011010101001010100000010100011001001000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out306[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out306, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100100010001100110011011101111011110011101011111011110101001001111101000111001101011100011110011101110011001101000001001000; 
out307 = 128'b10010110100001010111101101110001100110100000100010011011010111100110001000001100111001110000010011110011101010010100000100011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out307[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out307, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011010111100101100010100000101011111111100011101101100111100000100111111001111101101101100000101011111110101010011111100110; 
out308 = 128'b00111111001110100100011110010111100011110010111010000100110101111000101010001010010101110111100011010111001011000111101110101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out308[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out308, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001011010101110110000000000000101001100011101110001101111011011000000010010101111001100101100111110110100010110000101001011; 
out309 = 128'b11100011101101001100101000011110000110000111000110111101100100001111001111110110011001101101111011100000000000111010101110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out309[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out309, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101111110110100000011000001000110100000011101110100111110001001100100011011110001000111001001010010100001000110110100010110; 
out310 = 128'b10001000001001101101011011110011100011000101101101011000000000101011111010111010101000110110000111111001010000100101001100111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out310[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out310, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100010000000110100001001101011111111011001111111100100010110001011000011110000100100111110100000111010111000110001010011010; 
out311 = 128'b10000111010110010110000100010000011100010010010001101100101111000100111001110111111110100010000110001111101001011100100111011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out311[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out311, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111000111101001111000010001100000011110101101110110001001011110111011010011001000111000110111010111010001000100011010001111; 
out312 = 128'b01001111111011101011010000100101011010100110111110100110110111101000000001010110010110000110001011101001000001111011111011110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out312[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out312, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101000100110110111011011111011010101111011000000011110000001000111010011100111101111100001010111110011110100100010111010101; 
out313 = 128'b00010111010000100011000100001100001110001001101100010000101111011001100110100111110101101001001011011001001010001110011011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out313[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out313, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110110110001011001101000100000101111101000100010001111010011000010101101111000001110011000101010001010000001010111011110001; 
out314 = 128'b00110001000011001101111100000010111000000010110100110010100100001000010101110001111111111010111101001101000111111010010001101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out314[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out314, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000010001001111111010101100110010000110101100000101010011111010010110110001101100110001111111101011111111000110101100111100; 
out315 = 128'b00110101100001010110000111011000010110001110010001000010111010000110101011110101011011011010011001110001011001000001101001110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out315[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out315, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001000100000001101000011000000101100101110010101100000110110001000110101010010000100101110010100110110001111101111100100111; 
out316 = 128'b00011000100110100100101010010100101000111001100100110100111010111101100000100011101101110000111001100010100011010101110100101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out316[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out316, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100011010101011101111010011000010110000011110110010000010100111000001100010011110110011011011111000000010110101000100110110100; 
out317 = 128'b11110010101100011100110101101101101001000001000101100011111110100001011011011011011101111111000111000101001100011100110010001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out317[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out317, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001010101111000010100010000101100111111010000101001110011101111110001111011100000001110111101101000001000111110011100111001010; 
out318 = 128'b01101111001111111111001001100101011100100111011101001010001111011111000011010001101111111111000011000010111001111100101001111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out318[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out318, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100001001110000101100100011101001001011001010010000101111000011010001010000000000101111100010111011100111000100010001111100; 
out319 = 128'b01100100101111110011000010101101000100100010110011010001111001111000011110100011111000110010100111010000001000001010010000000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out319[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out319, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000010100010101001111000011000001101001000101101010010111101101101100110010010000000100001010111010010110010001101101101101; 
out320 = 128'b10101101111001101101111110011100010101101100111101110110100011101010000010101011110101011000110111110011100101000000001000111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out320[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out320, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110001000000100111110000100000100110101000111010010101010011101101111100000101000000010010010101101100000010111010000011101; 
out321 = 128'b01111111001011100101010001101111101100100101101001100100010110101100011111101101111101011010101010100000011110000001001011011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out321[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out321, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111100111110100111000100110011000001100100001010000000010111100000011100010111001010101100010010101011110111100000101000110; 
out322 = 128'b11001000100101000001010001101010111100100101011100010001000010100000110111001001101010010110011100010111001001100011001111011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out322[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out322, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001111011010010001011101010100010001001101100100100011011011010110001001111100100010011010111111011100010010111010110001011; 
out323 = 128'b11010011110000011110100010000111011100001011000110110001101010011010101110001011110000000001011010010101001010111001100100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out323[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out323, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110010110111111101101100111001001010000001110101111101111110111100001111101011011111001010111011101100010011010010001110010; 
out324 = 128'b01001101110110010001001110101110001010111000101101010101111110001111100110010101011111100101100100110101100010001000000100010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out324[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out324, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000111100101011111000100101010111111110000110000000011010000100100010111111001011100110101110010010000111011011011100001111000; 
out325 = 128'b11100010111001101111100000010111110011011000000111000110101101000000001011010001111011010101100111100110010110100011010111011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out325[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out325, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001010110000100111000000101001000101001000111110100100110000000001100111000110111110101111111011101111111000011110111110110; 
out326 = 128'b10111111000110001110010010100010111001100001011010011100100001011101000000010001010110011000010101110101000101110000110010000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out326[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out326, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001001110101100010000100110001100011011001111110110111100111011001000101110101100110111001001010011101001100101011010111100; 
out327 = 128'b11001000100101111100111011100000100101001111110101010111001000110010111111010010111111101101110101010100110100000011101101101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out327[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out327, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111011101111101111001001011101000101110111010111000010001100111001110100111011101000000011111101000001011010000101100001011; 
out328 = 128'b10111101101110010100111111110000001000101010101000101111101110111101101000011110000100110111110010001011101010111101000101111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out328[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out328, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001000010101011101100001011010101000010110000010011111010001100001000100010001100010010010010111011010101000101101100011001; 
out329 = 128'b10100010111101101111010001110010100101011001111111100111001101100001001100101010101100001001110001011101000011100011100100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out329[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out329, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011001010001110111100001111100011011000011110011001000110010110001111011001001101101101001011011001101100101111001100001100; 
out330 = 128'b11000010000100000101101010001011111101011111010011110101111011110011111010100111111011001010101100101101010111111010100111111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out330[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out330, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101100111111110101011100001010010010001100010111111101000111001010100010010001110111101110010101111011011100011000101001110; 
out331 = 128'b11000001010111100010001111011001011100001110111011110100000001100000111010101111000100011000011110100110010000010110110101101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out331[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out331, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011101110101110001110001111010101110111101100101110001111010010111011000011001011100000011110001111001001001101001000111101; 
out332 = 128'b00001111100111010110010111011101011001011001000011001101111010100100010111111101111000110100011110000101100001000010000001010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out332[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out332, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011101111010110010110011000111111011010111010000101100111101001100110110010110101011011000010100011101110111010010100001000; 
out333 = 128'b10110100011110010010101010110110100011000011111101000010101001001101110111010100011000111000011100001110001011011101000110101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out333[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out333, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000000110100011010110000100110000101010010010100000011111111000110001100100011011110011100000100011110011101111010100001101; 
out334 = 128'b11011100110000101100001101011110111110011110011101011101111001111011010000110100110011001000000100110111100100111000110001000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out334[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out334, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011011110010101100010001101110100011111110001101110000000111001111110110011011000001100000011010100111010001111011011100100; 
out335 = 128'b01010010110010000111111000110011100011111111110101000111001101000001110100110110101010011110001001100110101000110100010001101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out335[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out335, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101101101110001111000110001110001101000001010100110101110101011000001111000011101011011001101001001000100111100110000001110; 
out336 = 128'b00010101110110010101010111111000110011111001001110111100010000011101110100110101111000110011001011111110110000110000011111101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out336[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out336, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011110001110110110111101010111010111100011111110011010100111001001011110101000001101101101001010101010010111101011111011110; 
out337 = 128'b11111010110001110011011000000100111010010011101000000101101100100110110101100010101000111000010110011100010110010100101001000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out337[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out337, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110010000101011010000011001101111011011110100010000011111000000010001010101010010001101011101011000100001100001101001101101; 
out338 = 128'b00101110011100100111001000010000101110110110001101110001010010000101010100101110011011100101111001000110010010011010001110110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out338[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out338, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011010111111011001100001010110101001010100000000011011010110011010101000010000011000101111011001000001100110101000101001010; 
out339 = 128'b11010101001011010001001001101101110101000011011110110010010000110001101111100011011000010111111011100101000100101010010001101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out339[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out339, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110000111011101111111000111011001100110101110000101101101011100000110111010000011000101100011110010000010110010100001100000; 
out340 = 128'b01001100111101110011001000000000011100011010111110001111010010000010001110111010001101001100100000001011011101010000101011101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out340[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out340, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011000011110011111010011101110011101001101110010100111001101000010100001111010011010101010011111111101101111100101110111100; 
out341 = 128'b01110001110110111001010000111000100010010011100111001000011011010100000111111010011001000101000101000100111100001101011110111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out341[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out341, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110110000111001010011011011001111000100000010010000011010111100101111011100001000000001101110011100110000001000001110101001; 
out342 = 128'b10010100111000110101101111000011110011100110110100001001010000101110100111000100110110000110111101110100110000110101111001110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out342[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out342, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110001000000000110011111111000000000111010111010111010000111011101010010100001110110100101101011000111000011000011011110000; 
out343 = 128'b10010101001000001100000001100111111001001011110110001010110101011111010111000111110000000101100101001000110101000010001101111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out343[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out343, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111001101001010110000110100110111101101011011011101110010000110110110011100010100100011001110110111101010111111110001101101; 
out344 = 128'b11110100101011100011100111010000011001001001000111101110001011101001001000101111100101100000110000100101101001011111000111110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out344[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out344, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110000001011101101011001110000011100011100011010010110101010000011011011000111010101001000110010100110010100101000010100111110; 
out345 = 128'b10011111100000101010001000011011101110111010001101000000000111101101101001100010101001001000101001010001100100101011101001101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out345[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out345, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001001000101100100100110111010100001001000001111101010101110000000111000100010000101100001100010011110000010001100010111000; 
out346 = 128'b01000110010100111011000011100110100010000001101001001100001100110111110010000111110111010101011111000001010100100011000000011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out346[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out346, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001100001011100110111011111101000110001010000110110010100010111111100000001011010010001001111001100001011000011101001101011; 
out347 = 128'b10001001010001001101000100001001000110111000001010100111100001111101010111010011101111100101110100010100110000010000110100010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out347[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out347, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110101100100000101010110001000000111001110011100010110010100000111110101110001111001010110000110001110110000100000011111001; 
out348 = 128'b11001001010111110110011110000000001100110010000000010101110111101100111011101101100110001111010100100110011001110100000100011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out348[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out348, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111000111011101010111100001111111000000011001110010110000010100010100001110001001100111110111000101111101010001011100110011; 
out349 = 128'b01001011000111011110110101111101100010111000000011101000000100011111001101111010000000011100111111011011000010010101010100111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out349[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out349, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100110010100101001100000111100001000101011000010011001111001101111011101110001110101001000100001110101100100001001011001010; 
out350 = 128'b11001100100011100101010010011110001100111000001111011101110010000101000100000011100101000011101010111100001100000110100100011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out350[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out350, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110100000010011101111011010111010001100100111100101011101000001100011110100001001001100000001000111001000100010011101010001; 
out351 = 128'b01010001100001001100010110100111111110100000010101100000011000011100001100100110100101010001000011111101100110001001101011010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out351[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out351, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001001110001100010100110011101111011110100111111001101010010010101010110011110000100011111100101101110111100001101101000001; 
out352 = 128'b10111011111010110000000011101110011101010001100011001111111101111000101100101111010010001001011001110011000111010110110100101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out352[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out352, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110011101100100010111001001101011011101011111110110010100110101000110101110111100000010101111111010010100001011100100100111; 
out353 = 128'b01110110011010011001010010110010001010111010101001001011101001011000110110110010111101111100111000101111010111100101001000000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out353[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out353, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011100010000011011001000111000110000100011110100101011010010101011111000011100011011011101000110000001010111111010101001111; 
out354 = 128'b11110000110110111100110010000011001010001111010001100011010000110010011000000110110101101000111011101010010100000100110011100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out354[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out354, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011010000001011100001111100100101110010010011001000100011000100111101111010101100011010110000011101100010111111100110011010; 
out355 = 128'b10111101001111000100100101110101001011011100001011110001111000100101000010001011100000000010010000110010001111110001011100110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out355[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out355, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101010100011111101010001100111011100101010111010000110000000100100011000011101101001000110101011110000110101011111011011001; 
out356 = 128'b11000100101010111111100011001110111111110111100001001101000100010110011001000010111110000001111001100011100000110011110100001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out356[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out356, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111101010001111110010010110101001010111111110110111001101100010001101100001110101101000001001010110101100011011110100101111011; 
out357 = 128'b01010111010111000010010010001101011010101001101110111001010101010010000100100001011010110011110011101011000101100110100011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out357[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out357, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111110010100110001011111101110011100010111010110011110000110101000011000011111111110101000010101110000110111101110111010010101; 
out358 = 128'b00011001011001000110001100000111101101011001110010010000111110011011110000110101001001000100001000000001111100001010110011010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out358[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out358, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111011011001101011011001101010101100111001100011110100000000101100010111111001110001111001111000001101111011010110011111000; 
out359 = 128'b00001001001111011111110001010001100110100010011001010000011001011101010100011000010110110010001000111010100011011100000001010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out359[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out359, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111010001110100100010100111110001010011101100011101100011011110001110100011101111101110111010000100011010011001100110011111; 
out360 = 128'b11011000100000000010010001011010010000100101011111001111010101010111100111100110110101000010101110000100010001000110010110000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out360[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out360, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100001011111111110111001010010101111101000111011101010101100100101101101001000000111000010110100010111001110010111001001111; 
out361 = 128'b01011100010100100010100000011000011000010110011010010101011110111010110010110010111010111010001111111000011001100010110001111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out361[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out361, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110011011100111010010011011011100000111010001111111001111000110110001001010011101111000000011011110010111000111110011000101; 
out362 = 128'b11000100011000100100000101110011110100111011011010111101111101110111000011001001001110110111010111100110010100111100100000010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out362[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out362, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110000110100001111000011100100110101011100001111011110100000000101101010011001011111110110010000110100001001110110001011111; 
out363 = 128'b11110100010110000101111100001010001011101000010010001100110001011101000111001110110001000011110011100101000011010011111100001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out363[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out363, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110001110101011101011100001011001000010000100001111110101000000010010100100110011000101011100001011000010100111000101010111; 
out364 = 128'b11100101000011110100001011000011001111011000000110011110111011001010100100011110111100101101001001100101001111100100111000010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out364[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out364, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110101111111110000101101010101111111000101010110010010100111010110100001100000010011001101101100000101000010000100001100000; 
out365 = 128'b10001100010111000100100010000010111110011011000111010000101111010000110111101111001000011110111101010011111001101011000100000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out365[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out365, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001111011000010011010010010001000111000100011010100001100000000000110100101000100001111000010001010110001010111110010010111000; 
out366 = 128'b11000101001010010010011111001011010100111001001101100100011110001000101001001001111111000011000010001100000110010101110011001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out366[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out366, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111110101011101100101111000101111001010010101001000101011101110011100110011010011011010010010100101010011001101111111100101; 
out367 = 128'b01101101000001101110010101001110001011001110101010010101101000000101010000000111111101100000010101101101011111011011010010011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out367[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out367, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101010001111110101110011111010000101110100011110110100000011100101110111011011000010000010001001100101100111000010101000110; 
out368 = 128'b10010100110011011101110100100000101001100111100001111110011101000000011011100010010001101010110001101111101111100111111111001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out368[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out368, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011100110101011110010001011000010010101000011011110100001111001011000000101010000000111001100000010110101001110010101101101111; 
out369 = 128'b00011000111100011010101011110001010111110100011011110001110101110101001111010100010111111001111101010111001011000001101111100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out369[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out369, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110110110100001111001100110001111010110101011110010101110110100010000100100110000001011010010011101001100011111000110101001; 
out370 = 128'b00101100001011101011110001101100010001001010100001111000010011110010111110000011010001111000000100011011101100011111001000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out370[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out370, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001100110110001011110100111001010011101011100011010111000100010111001111011110111101011011110100011101110101001111001101101; 
out371 = 128'b10011000011110011111001111100011010011101111100011111011110110011101010110011011110101001000110011101110010001011101000011010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out371[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out371, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110100001111011011101111110000101100010100101100011100010011000001011011001011101101100001011111110111000110111100110101100; 
out372 = 128'b11101010111101110111010001000010100101001000101101011001101010111011011000101010001101010010110010001110001001010010111101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out372[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out372, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101100110001000011100101010010000111100101100011101100000101110110110110100011000100011001010000010001100001011101110011110; 
out373 = 128'b00011001101111001101101111100101011001101101000111011010110101011100101110000011011100000111001011000011010111111001001001000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out373[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out373, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100111111001101110111101001101100001010100110100000110110100101110111110111100011000110100010000111111011000001000100010001; 
out374 = 128'b00111111000011001000101110111111111110111101001101010010101111100100001111100100101000010010111110100111101011011101110010010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out374[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out374, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010110001000101101100101100011010110001001011010011010111001001101011000001101111100100000111011110001000001100010010100010; 
out375 = 128'b01111011011110110101000000101011101100001101010110011000101011101100001110001010111110011000101101100111111011110001000111001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out375[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out375, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000011001000100001101001101100111000001001101101100101111111100111011000101001001000010111111010010010011110100010111000000; 
out376 = 128'b11111100000010110110101001011001101001011101100110111010100110100010000000010001100010101110110111111110011001110000111100000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out376[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out376, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101011100111011111100101000110101101111111111000110011010100000111101001000011001100010111000010000011101011101100110100000; 
out377 = 128'b00011011111011011100100111100111010100110000011010100110010111001100111011100011111010100111001101001010001010010000011110001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out377[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out377, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111011101101110011011110101110111001111101100001111000111001001011101100011100010101101001110101011000100000111110101001010; 
out378 = 128'b11001011010011111111000100000111100111111001100111111011000111101101100110001110111011011101100100000011000100001101011001010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out378[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out378, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010100011000101000001100110011111000111111100011011111111010100000001011111100010011010100101110100001100011100100001111011; 
out379 = 128'b01001011111110110101000001111000011110010011001111101001100011011101101011001001000110101100101101000001000010111101010011111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out379[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out379, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110000011100001000100110101010111110010010110000111000101110001001010110110100101111100000010000101011000111000010100001010; 
out380 = 128'b01001111101100111010000011100110100000001101000101011000011111101000001111000111101010110110110010110010111001110111101100100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out380[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out380, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101100010101110000111000101111110001101010101011111010100101011001010011111001111101111110011000110110001011011101100010000; 
out381 = 128'b10111101100111010001101000111000010011110101100110001100100100100110010011101101010000110000010011111000010011011110100011101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out381[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out381, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001001000111100100000011101010010100011001011101111111011010101000110001100000000001000110111110100000101000000111000000101100; 
out382 = 128'b10101010101101100100010001100010110111100101011010100100011110001100001000100101110100001011000110011100100100101010110001100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out382[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out382, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001101011101010001010110111001000011100110001010001100111111110110001001011100010111001110101111011001001000001000100110110; 
out383 = 128'b10111111010011111100001101001010001010100001010001000110111110000101101100011000100100110111010011011011000001111010101001000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out383[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out383, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110011111011010110010010100000001101110010001000011011001101101010101101011101100101110101101111010001111010111000111100111; 
out384 = 128'b11010101100111010110000110010000011011101111010101111001011111001101101100100101111000011111010111011010110110100001011011101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out384[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out384, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111101100100100001001000101100101011101111111000000100011010110100111001101011011010100010111101100110111101111100011101000; 
out385 = 128'b01010000111100110100101010011100000000010010011101111111110100110000100101001100011010000111101011011110010010010001000101111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out385[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out385, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101010001010000110000011111001101110000101001000001001011000110011001110100000110110011111111110011110110011010000101110101; 
out386 = 128'b00110010111100101000100100110101010011011111000100011001001111011011010001101011100101011101001101001101101110001111110000000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out386[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out386, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011101110000111111010001010011111000001000010101000011001100011100011101011101001010100100101010010110000101111001000100110; 
out387 = 128'b01111011000011010000110001010011110101011010001000111101010101010001001110110110000001110010110110110010010110010110111011110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out387[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out387, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110100000001011010111001000000000101010110100110010100000111111111110110000010011100101001100111010010010000011011001000011; 
out388 = 128'b00101001101011011000011011111111000110111001110001010000000100011001111001001011001110000000100001110000001001001101110101101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out388[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out388, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100111010000101100111010001101000011001101011110100100110110100001110101001100001010010011111011000010001000101110101100000; 
out389 = 128'b10000000001111001111110010100010010100000111010001011000000101010001111011110100010010010110011000000000000100100100001011111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out389[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out389, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001000000011101010011001010001100101110001001011010010110000111011100011101111001000011010010011001100110011010000011010001; 
out390 = 128'b01010100011010111110010101010110110010111100011010111110010001011000111101011000011101010000111101100010001001111010000000100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out390[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out390, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101001010000011000010101111101010101011010001101111100001000011011111100101111100110110011000101001101001010010101001000100; 
out391 = 128'b10010000110111110000101011000110110010010100001100100111000000010110011101011000000111111110100111001100110100111011011001101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out391[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out391, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001010000100000100000010000010101101110100100100011010111101110101110000100111110110001111101010101001000111001001010101111; 
out392 = 128'b11110001101010110101000000000010001100010000111001101111001111101101001100010100011011111011000010011010100110101010011000101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out392[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out392, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010110001000101110100110010111100010010000110010000010101000001011010110101110110010000100010000011110111010111011110000000; 
out393 = 128'b00000110011101100001001010000010000101010011001110001111010101011110010001010000110111010010010011110011011101010010110101001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out393[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out393, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100101100110010011110111111000111100100011001110111100011100111011110111111111111100101110100011011101001110000000000000010010; 
out394 = 128'b00001010000110010011001010010000011111011101111010100101111011110011010011000010100101111000011001101111110011101001010111111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out394[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out394, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101001001000011010001011101011111110011001001000001110000011110111010101010001000001111111001110001101100100100011100111100; 
out395 = 128'b00001011111001101101011100001011110101011101110011100011110000111010010011011001011110000011001011110111111111111010111001010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out395[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out395, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110000101100011110110101011100101001111010011010101001111011111001001101111111000101001001010100111101100001110010111111110001; 
out396 = 128'b11001101001100101110001011001100111011011010110100011001100000001011110100010011011101110000000110011110011011011010101000111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out396[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out396, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111100001001010000001001111000010101011100110001000100000100011011101110001100000111001101101011111101110100001101100010010; 
out397 = 128'b01100100010111101010101100011101111110000110011111010110000011101010010110100010101001000000000011010100000000111100100110111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out397[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out397, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111111001100100000011011111111110001000101001111101001001101111010111101011101000000111001011110001000011000110001111000000; 
out398 = 128'b00011001110111100110010101011000110111000110010010000000001110011010011100000010111010111001111110110100011101110101000001000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out398[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out398, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001100001101100111011110010101100011100000011111111011011111010101100111100000011010001000111110111010001111000111001010011; 
out399 = 128'b10000011001101101110001010000101111100010011011110011110011011101100101101110100111001110000010011010111010010101000011000000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out399[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out399, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100100100100100010110100101001100100100111100100010100101101001001101110110100010101101100001100000111100110010111100001001; 
out400 = 128'b10100001111010101111101101001011110011111011101101000010100100010100010111011101011011101000110001111011101111101011011011111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out400[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out400, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111101111010000110011111111000001000000010101100000110010001000101110001010100100010001011110010011110101110011100110101011111; 
out401 = 128'b11101010111011111110111100110111011011001101101011100111010000111010100110100111100011001111010111111000110011100000010000001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out401[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out401, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001101111010110010011110110101100001111010000110111100100011111010111110011011001110000100000001100110000001000000101011001; 
out402 = 128'b00011101011001111111101011001101001000101000111101001000110001111110000001110011011001110110011000001101011010000000111000101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out402[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out402, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111110010111010100110010000010111101110100100010111100000100000001011011100110000101001111111011100001111000000111001100010; 
out403 = 128'b11010010111101000010001111011101110001011010101100111100110100000011101000100001101011000000010011011101110011010100101010100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out403[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out403, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111000111110010000011110010001101001111000011100101011000100100101101101011010110100110001010001110000100001000110001111000; 
out404 = 128'b10100100001100100110111001001100111001110011011011011111100011110100110010001001001111001110000011001111011110011001110011010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out404[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out404, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011101110100100111000010010111001111010001100010001000000001010111101111000100010101111000000111101101001011101000011011110; 
out405 = 128'b00010010110100110111000001011101001000110010111110010111101001011001101101101010001110101101110010000100000011000010110100010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out405[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out405, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011011101111110101010001101001011010010101110110101111011001010011000111110111000000010100000000100110101100011010111000011; 
out406 = 128'b11100100010111010111100111110011000001001111001101101110110110011010001001010010100011000101100111011111100011011001010010010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out406[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out406, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100010011101011001110010011011111100111111001111001101101110101111010111010010100011100010010110010000011111010100011010101011; 
out407 = 128'b10001110101011011011001101001000011110000110110111011011011010011111001111101101010010010100011000011000110111011011000001100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out407[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out407, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100011101001011110101011111001001110101101011000101111000101111101011010010110011000010010110110010011010001001010000001001; 
out408 = 128'b10001000011010110011111000110001110111101000001011111100001101101000000100111001001001010001111101001011100101111100010101110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out408[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out408, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111111011111110001101010011010111000001010101010100001110101110101011011011101011001111111101011110011100011001101011010110; 
out409 = 128'b10010110011111110100000110001001101100001011011010111001010000110001011110011011110010000100010000010110010111001001111110011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out409[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out409, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000010001011111001001100001000111110101000100010000110001000000010010000000111100001100110010011001010110010000110011101011; 
out410 = 128'b00011110101010101000100010011100011111111010000110101000110111011011011010100000101011001000110011100110010000011111100000101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out410[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out410, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001011100100100101100100010101000000101110011111100100101001100010101010011010100110111011011111100111111110011110101101100; 
out411 = 128'b11110110011110001010100111100010100101100110000100011011011001000101011001100011011100011001111010010000101101100101000000010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out411[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out411, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110110101011100011000010110001101001101010011100100111101100110000110100100010001101101110011010001001110100010100111100110; 
out412 = 128'b11001101110100110110010110010101000011001100101101001000111001011101001111110010100000011101010010001010101010110001110100101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out412[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out412, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000011101010000001011110010110101110111101000100011111101011011010000101000110100010000101000011111001100010010001100110111; 
out413 = 128'b11100011101001010000010001110010010110100000000101100110101001101000000101100011000101001010100101011001001110000100111101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out413[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out413, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110000100101111100111000111111001011101101111110010001111010111101100011011011000100000001100001010111110011110100101001101; 
out414 = 128'b10000111101010001011101000101010110010001111110010010010010011110110010010000110101101001111110101110000101011001110110110001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out414[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out414, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001101001101001100100000010000001011100001011001000010100100000110100000100000011001010000110101101100111111111010111111001111; 
out415 = 128'b10111111110111011110011000000100110110101010010100001010000011011000011100111100100110001111100111110001101010111101000001010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out415[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out415, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001110110100001100101001011010100101101011000111100010010011011000110001011111110001011110001001101110000100001111010111111; 
out416 = 128'b01001011101000001001001111001111010110111110000101100110001111100000100000110010100000011100101100010001001101001010011000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out416[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out416, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100101111101000101111011000010101001101010000110000010111101111010000010010010110011001011001000100111001000001101111011010; 
out417 = 128'b11101100010100110101110100000010101011101001110011011011101100000000010011001011001100011100010111011001000010101100000011001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out417[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out417, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001110101000001000000100011110010001111010100001110011101100001111110111100110000110100000101000010001101101110100001111000100; 
out418 = 128'b11110101011011011100100111110101110011011100110000011101110111110011111110101110001011011011111101010000100011110101001111101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out418[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out418, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001010100010010001100010010111110111000010011000001011011111001010110100010110110101110100101010110001110101001111110100100; 
out419 = 128'b01111110110010101111000010111101101011101101000000000010101010000001101100000111001110001111010010000011101110111110001111100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out419[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out419, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000011111100001011101111000110010110111001000010010000111111110011110000011010001100111001100001001111100011011110010111110; 
out420 = 128'b01001011101010100001101110001010101001101001010010110101011101000000011010100000101110110110000110111100010011010110000001111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out420[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out420, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011101110011110010100110110011110100110010001100100010100101100010100110000111001010111110011000000000111101001111000100111; 
out421 = 128'b11110001000010101000000100110011011111111101111111111101011011001110010111010000001101100111001000110101100000111000011011001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out421[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out421, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111111001101101100001100101010011001001000000110010111010011111100011001101010000111000111010011011110001110110101110011111; 
out422 = 128'b11110100000101101000111110111100011100000111101110101110000111000111010010010110100011101111111110110011101010101110010110100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out422[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out422, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000001101100010000100001101000111110110011101010011010110100110011100110101101100001001000110011010011010101010101000100001; 
out423 = 128'b10111010001011101111001011101110110111010010110011110101000101010111010011010010001000110101100000010100101001010100100001100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out423[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out423, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111000100111000001111100011101100100010011000110101010001110000011000001000000110000000000111001001111100000100010010100011; 
out424 = 128'b01100000010000011000110111001101010101011100000110100111000101101010001111001010000010111100100010000000011101000001111110010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out424[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out424, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000100101101011111111101100001101001000010000101000001011111001000110000110111001000110001011111110001011111010111111110110000; 
out425 = 128'b11110110000101010101100010111101000000010001000010100000101010011000000111000000000111101111010001010000010111100101100001100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out425[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out425, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100000101000010001101111101110111101100000010010101000001100010101101001100100011000010011100110101011010111101001100111001011; 
out426 = 128'b10000110110111000011011110000100111110000000001100110010000101101110011100000100010100010000111000100010110110100100101001010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out426[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out426, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001010110010011101000010110110101100001010000101010110010101100011011010000000111000110100010100000000110111001101011100111; 
out427 = 128'b11010110000000010110101001111111000101000001111100000110110100111101111111010111110010000000110100011111110100111111011010010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out427[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out427, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010000010101011110111110110110000110011010100011100101011111000001011000111110101111111110001111101100111111010101100011001; 
out428 = 128'b01010100011001100001000101111110001001101000011001100100011111010111011110101110011100101111110001000000111100000010000000010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out428[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out428, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000100111010100111111010011100100100011111000001110001100000000010000111100100110100101011101110010010110010001110011110110; 
out429 = 128'b00110010111001101110001001111111000000100111100111010110001101111111101011011100011110011100110011101010010001101111100010000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out429[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out429, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100000100101010011011010110011011011101011011000010111000011101011100111101110111110010101111101100100001101101001101100111110; 
out430 = 128'b00101110101101000110010011010110010100000000010110010111101111011000000101000100001100101001101110000100011000011000100001001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out430[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out430, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100110010010110100001100010111110101000100000011110110001001001100111010101101001011100000111110000111010010111011110100011; 
out431 = 128'b01111010000001011110010001101010101101101000111010010101001000001000110111011010001011010001011110100101100101100000100110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out431[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out431, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111111101100111010010000111000000011011011100101010110010101001010001101000001100101111110111101010000110111111000111110001; 
out432 = 128'b11101001101101001011101010011101100101011010001010100011011010111001001110000000011010101100000111111001000001010000110111100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out432[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out432, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100011110100100100110000101111000110010011101110010100101011101000110100111100010101000011001101101000101010000010101001111; 
out433 = 128'b10111110110101011011111100110100110001011111111111011110111011011100100010000010010000111110011011100001000100101101100000111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out433[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out433, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101110010111001001100100001001100110111010110011111110101101110011100011000111101110100010101111000110111101110011010111011; 
out434 = 128'b00111001001110100101111111100000010010100111110111100010000100100111010010010101010010100110111111101011001011110010110001010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out434[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out434, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101001000001001101010010001111111111010101110010110110001101000010000010001010001111011010101101000011111010000001110100011; 
out435 = 128'b10010011011101010100110100001010110000111001011111100011101010000011111001010000100111000011101101110000110110101011100110101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out435[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out435, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010001000100000001110001011101100110010001111011001101010011100011000001101101001000010000101001010001010111011100010111100111; 
out436 = 128'b00110010100001010010110110001101101110100101001010011000010110111101100011111111101000010100010011111100110100100011011010010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out436[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out436, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001001001111101010110111110111000101100011101011111111000001010001000001110100010111011100010011111110110100010001100011110; 
out437 = 128'b11010011111001010011001100011010010111010100011000100111101101111001110101000000110101100101011010111100010011101101111110001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out437[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out437, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110000111100100110100111101000000101000100001100001011011101110110100111011010000011011011001010110101101010000110111100000; 
out438 = 128'b11111100100111010000101000101010100001111101001111101000110000100000011111110000100110110101000000001100001111000000011001001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out438[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out438, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001111101110000101110010000101110111010101000110110110010000011010011100000111001110100000111100011110001000001011110010000; 
out439 = 128'b11101101011111001100111110100000000000010101100101001101110000110000001000010001100010001011001100000001000001010001101010011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out439[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out439, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110101000001100000110110011111110011011001001001000101101101111010000111110010000011101001110001101011011101100011011000100; 
out440 = 128'b10101000010110010000110010001000110110110110110000010100101001111111101011011001101000010000001100011111101000001010011011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out440[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out440, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110001011001111000110100000010100011001111000011101111011000100000000101110010110100101110111111101000000100010100011010011; 
out441 = 128'b11100100011111001111000110010010001100110010110110111010101111000101010100110110110010111001100011110100100000001110000011111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out441[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out441, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111000101011101111001010100010110100110111011000001011111100100011100111111000000011110100001010110111010001001011101010100; 
out442 = 128'b11000010111011010001000110000010100001110101011001000101010000000100110110111101101101011111001111010111101101001010110101010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out442[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out442, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100111100101001111110110001000111101110011100110110010010010001111111001000100110010110001101100100011001110011101000010110; 
out443 = 128'b01111011111111101101110000101000111011011010110011001110001100100011110100011001100000000000000101110000011101110101101011000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out443[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out443, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100100100000110101101101111001110100101001001110111111000101101010110010010010111110100011001001111000100110111000001111001; 
out444 = 128'b01001100011110001110110010111010110011110110011100100100010001000111100000111011110000101110110100111011100010111110001111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out444[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out444, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101111101111000111111001101010000011111010010000111011011110000010000101011000100110110010011100110010111001111010010010010; 
out445 = 128'b00110110110110011110100111100101011000110011000110001000011111010010001010000000110101000010111000000101100001011100100000101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out445[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out445, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010111111000000100001110101011100000111000111000101000001010000001110001010101011101101010100110000101011101111010000101010; 
out446 = 128'b10011001110101000101001000011110010100001011100000010101110111111100101100101100111110100010101100101001011010110011101111010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out446[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out446, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100000101101010100011011100000011111010001011000000001000101110111100111000010001001001000000100110100000110110010000110001; 
out447 = 128'b00011111010010010000011010111111010000000101101101001111010010111100010001001000100111110001100110111110010001001100101100111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out447[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out447, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001100100011110111110110010010000111111111011110001101010010000010000011100111001110000001011111101111101010100100011101110; 
out448 = 128'b01001111000100111100101100011100000011111001110001100111010010010000000100111101101000011110010000111101100010000011111101101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out448[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out448, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111100011100101010110100010111000100000101010001111011111001110011010000001011001111110100001100100101010000100110001011000; 
out449 = 128'b00110001111001011101111001110000100000111010101101000110010101010110000001010101101110010101100000011101100000100011100010010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out449[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out449, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110111010010011011001111100110111011110000100100100100110011111100011001000001000110101001111000110101001010011000000101010; 
out450 = 128'b10101101100111001110001101000111000100111001110110011000110001010100010001010000000111100000111110011101010101100001001111001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out450[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out450, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111111010101101000001111111110100000000000010011110000110100001100011111100111011101011101110100011110011100000011010001011; 
out451 = 128'b00000100111110110011011100111000000111110010100000001110111111011010100000100001010011111111011100010101101000101000100101010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out451[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out451, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001000101101110101111000010111101111011010111101010100001000101101011101111111110000001111100001001100011101010111110001100011; 
out452 = 128'b10001110000010110111010101001011000001100110111100011000111000000110001101000011000010011000110010000101000011101001001010011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out452[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out452, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110010101111001111101100111001110110110100111010100111010110000101011110100010010011101101000100011011110001100011011111111; 
out453 = 128'b01111111011000111110111010000101110000001010100110101000110010001100110100000110011100000000101000011011010001000001101000001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out453[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out453, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011101111000110011101010100011110000010000111011011001111000011100000010111000010010011110100110101000110111010000011000101; 
out454 = 128'b01011001011111101101111111100010101100001000001010001001101000101111100011000110001100100111001001000110000111011011001001100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out454[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out454, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111111000011110000101111000011010000111001011111001001001101110010000001010011010010101101101010001010101001110100111101011; 
out455 = 128'b10110001100000010100100000111010110100110000001110011010001100011101011101010111011000000010010100111010001101101111001101001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out455[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out455, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000101010001010000011010101111101001001000010111111001011001100101010100100110010001010000100110001111000101011011101011011; 
out456 = 128'b00100010101010000111111111110101001011101110001111100000010101100001000010101110011001101111110101100100010001111100111101110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out456[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out456, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101100100100001111010110101011010111001100000100100011101100100100011111110000110110110101100010111011101010000000000010001; 
out457 = 128'b00101001000111100101010001101010100110010001000100001111011110010111000100011011010011010100000111100000010001110000101100110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out457[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out457, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100010111011110111001110010011111100101000111000010110101100011101001011000101001011000010111111110000010011101010100011010; 
out458 = 128'b00100001010110100110110100011100100101101011001100011100110011000001011100011100101110111000100011111001010101011111011110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out458[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out458, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110010001101001100010101101011010011111100011100011000111000111111101110111001011101001101011011000000000111011001010011110; 
out459 = 128'b01101011000111111011011100111101000011110111110110100100011110101000000110000000000101011101100111010100011000010000100110100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out459[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out459, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111101111000100101101001100110110111101001000000110110100010111100110100111000100111000010010101100100110001111110011000000; 
out460 = 128'b00101011110010110101011111111011011011110001100001011001011011110101010111011011001100010100010001111010110010011100101110101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out460[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out460, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001000001011011110011100010110010110101111101000100101110001000101010011100010011110010100000110001011011010000000101111111; 
out461 = 128'b01101110000111101010101111011000000111000011000010101010011001001100011101011010011110111001111101001001011101111100011111111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out461[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out461, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000011100001110101000100110011001111001001111100001010110101010010000110110100010101010000101011100101011100000100010001101; 
out462 = 128'b00011011110100010010110011000011000101011101011010011011101111111010101101010100101000000111111100010001100011010101010101100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out462[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out462, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001111100000111111001000000011100110101101011110100000111001100000001001100000010010010101000110000011011011111110001010111; 
out463 = 128'b10010111101101001110110011010110111111011110010110010000010100100101101010100100111011011100100101100110001001110001100111001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out463[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out463, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001101111110100111111010001100010111101101001101010110101110110011111000110100111001100011010010111100110111010101110010111; 
out464 = 128'b00010110010000101001011000010110101000001000111010010011000000100110011010001001100010001010011110100011000110011010110110110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out464[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out464, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100111111000100011110010011100001010011100100111110101111110011010001100111000110000101110100011010010001010110001111001101; 
out465 = 128'b01010010011110111010111011000100100110101100001111110000111011101100100111101101010001000001010000110001010101100011111000101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out465[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out465, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100011000011011001111111001101000000010111011111011111010010101110111011000011001111100000000100100100011101111001011101100111; 
out466 = 128'b00000100111011010011000011101110101011000000111111000101101110011101000110111101000100011001010100011000100110111011010100100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out466[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out466, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010010111111111000001011000111111111100011110010011111010110010000000001000010110110110000011000101000100101001111010000011; 
out467 = 128'b11111101100010010100000011101011111000000000101010100000011001000111011111101101100101100101011001010110011110101000010110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out467[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out467, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111001010100011001010000001100111110001110101000110110000010111101111110100011000001000110110111010111111110110111011101010100; 
out468 = 128'b11101110001101101101000010011000111110001111011101101001101000001010110001111011011111111101111111101100111100110101100110101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out468[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out468, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111111000001001001011010001010110011100110101101110110100111010100111000100100111010111011100110011000000001010010101001101; 
out469 = 128'b01101010101010101110111101010110100101011101000110100011111111111010110000000001100111110100000000010110010010111011101110011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out469[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out469, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010100100010101111101001000101000101000011101110111101111010110010101100001101101111011111000101100111100011001101010101100; 
out470 = 128'b10100001110110101101011000000000111011011000000010001000010100010001001110010110011011110011111111001011100110011111111000100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out470[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out470, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011101110100110000011001001001001100100010010010100111001011101001011110001010110110101011101110011110001101010100000101111; 
out471 = 128'b10001111001011000111011010100001011001110011001000100011011001000110110000100001101110100011000111011010101011110111110110011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out471[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out471, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001100100110010001000100101110010101011110100111001010111100110100101000100101000100000110001110110000000110100011100011101; 
out472 = 128'b10111011001010000011001101110001100100101111101010001110011011010101000100000111000001100101011000010010101110111111110001001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out472[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out472, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010100111011100100001100111100010010100001001111100101001011011010011111101000010110110011010100000010111101110110100001111; 
out473 = 128'b00111010101010100001101000110100111010101111010001100001100110111110011110111000111101111001010010011110110010110011101001011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out473[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out473, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010011000011100100000101001110011111011010111110101001101101101110110001110010011010011010000011010011101000011110100111011; 
out474 = 128'b01111001110001100111100111100110101111001110100001100111101010011101101011001101100110010011000001110111000111000011000010011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out474[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out474, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010110110110001000110000110000010101110001100110011101101100010111001010011010100011000011001011100111111011010100111101011; 
out475 = 128'b10010000001010001011011101101110110001000101001001011110001010111011110000011100001010011111011010001000010101001011101011110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out475[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out475, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000000110010001111101001000110011011001001101000101011111010100001111110001000010101011101100111010011100110001011000011110; 
out476 = 128'b11000011110110000111010101110011111010100101100010000001001101110110010010101001001110110110010111000001111011100010010111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out476[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out476, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001010110001000000111000001001100110011111000111101011101000000111001111001000011100001011010110100001011001001100110000101; 
out477 = 128'b10110011111011111110011000010010100001100001110110000011110001110010001000011001101011100010010000001100001111010101001001100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out477[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out477, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111101110000001001010110100110100100111001010110101001110111100111000011101110101110100010110110111000111001010000100101000; 
out478 = 128'b11010111011111011111101001011111110110001110001101100011010101100110000100000111101000110100101011111000110000111010100111111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out478[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out478, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010010011101000111000101000111111001011000111001011110001100010010001000001010000000011010001001000111011000110001110111000011; 
out479 = 128'b00100101000010000000000100011111001100101110001010011000001000111110111101111000011100100101010100110100111010100001111000110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out479[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out479, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011100010101001111111011011100100110110000010010000011111001010010100001001111101011100110110100100110111011000010010000001; 
out480 = 128'b11001000000001001011001111000011110100011110000010010101100001010001100011101111101000110100001101011010010111110010110000000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out480[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out480, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011100101100000001001011100011010111011001001101010001000000000010010001111001110101000010010001110111101101001010001101001; 
out481 = 128'b01000110100111101011001001111000111111100001010101101100010100111110000000011101010011111101010000110100011011111000110000011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out481[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out481, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100001010110101011101011110001111111110010111111111000111000100010101101011000101110000111001010100110101100110110010110101; 
out482 = 128'b01110011111001111100111000111011110101010010111000000010010100110111010010000011010010110001111011000000011010010000111000111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out482[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out482, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100111111000000100011100101000110010011110000111101111000010111101010010000001001001111001000111000011000001101001001100110; 
out483 = 128'b01100011110111010100101000101100011110100111011001111001011000110110011101011100110111001000101110100011110010000111010011111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out483[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out483, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100111000010011111100000010011111101011011001000010010111011101001100110110101110101001000110011100001000011100110010000101; 
out484 = 128'b11000000001110000000001110101001011011110111000010101010100111001101011101111001100101010101000011110100110111001110101001001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out484[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out484, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110001101010100011010100110011000100011001111010011100100110001011101010010001011101010101000110101011011001110011001011001; 
out485 = 128'b00111101101001110000011110001111101000000010111110100111010101110111001101010001001001101010101110000001111001101010111101010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out485[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out485, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100110011011111111011011011100111110011010011101000001010011011001110011100111101100110110001000001110000111110011100010101; 
out486 = 128'b10010110100110011101100011000110010000111011101000000110011110011101000010000100010100011111011101100011101011101001011001010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out486[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out486, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101011110100010010100100001100111101101101001001111000101111010111111100111111111011010101010001000000011011110010100001010; 
out487 = 128'b00101011101100000010101000000111001010011111111111011101000111001100010000111001110001101110010000011101100001110101111101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out487[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out487, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101010100100001111101111001001001000011010100000100011100011001111100001000101100100001010010111100100000000101000100100101; 
out488 = 128'b11000110100110001001010010010010001001110101101011011011110010011100111011010111011001011010010010110001000000010001001111010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out488[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out488, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101010011110100101101011101011100010001000011001001101101110100100110001001100010001010101110101100011011101001111101001010111; 
out489 = 128'b10101101001001000110000100010010011101110111010010110000001011011010110010010010000010111111001101000100011111000000000011110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out489[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out489, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110000100111111110110110011110101001011011100011011011000101110110000101001111001011010111111001111000010101110100100111000; 
out490 = 128'b10010110010110100010001100101000011110111001001001000111110110100101001100001111010110011001100000110001010110001010011110011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out490[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out490, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110111100110010100010111001101010011110100001101111100000001010010001110111010100011100000100110001001000000011101001011010; 
out491 = 128'b10001000110010011011011010011100001000110010111010000000100100000010101010111101011011100111101100000101100111010110000001011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out491[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out491, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110010101001011001010000011110011110100010011011010011111100110010001000001110000010010001101011111010010000000101010001000; 
out492 = 128'b10100100110001100101010101111101001101111011011000100110011010001101111001110101010010110010001001010001001010111100001011000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out492[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out492, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111011000110001001000011101001001110100010000000000000001111001000010110010000111001011011101111111000010100111100010011011; 
out493 = 128'b10100000111110001110011111010011010000111101101011100110010101100100000011001110110000010000001010010110011011000111001010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out493[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out493, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001000111000100100110001100100000101001011110101000001010010100110000000111001010011000100000011101000100101011100110000000; 
out494 = 128'b11011100010110010110111100110111011011001101000110111100001100110000010011111001011000110110010001010110110001010101001011000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out494[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out494, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111000111100110101110000001111111110110111100110000110011100011010110010100111111001001011111110110010101011011001010101101110; 
out495 = 128'b01100110000011101111101111001111000010100101011011111010010100000011000100001011001010111100110010001110111000000011011001100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out495[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out495, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101010000101000010001000111110001100000011111100010111010010011010000000111100101011001000010011011111000111011110101000111; 
out496 = 128'b00010100111011010100001110100011010000011110001111001111110011101011010100110010100001111001010001101100101111100011001011010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out496[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out496, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101111011111011000101100000001110111110100001110011000001011000100001101111001111100000001000101001010100111000000111011010; 
out497 = 128'b11011000111111110101101000000100111000111101010010101110110101011010110111101100000010100111110010100101100100010000011101000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out497[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out497, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000111010100001100010000111001000101001101101110110011011000010101111101001000000101100110000101111101010000010001110111001; 
out498 = 128'b00011110010101001010011110111001111101011100010110101001001011011000101101110110000011001011100011110110001010001111110110001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out498[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out498, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100110001001001100000111111111101001000111001100110001000101000111011100100110110101011011000101000000101000010010001110100; 
out499 = 128'b00100100000000100010011101001110111110011010101101111111101111101111110110010100110110101101000110010100100100001111000100111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out499[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out499, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111100010100111110000101011100011001110001111001110011001011011011101110011110001111010100110010111010001110000011011101001; 
out500 = 128'b10100000010010100011011101011011111111010111000000100111110011000011001111010010010101111011001001101100010110111101100010111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out500[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out500, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110000000100011100101110010001001010100110000010010111111010111000100010011000101111010001010010001000001101100101001000000; 
out501 = 128'b00010110000010001011110110110100100110111111111011110001101010111010111101010011011001100011110001000011110001100100111001111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out501[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out501, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000011100001011111101010011101100010010010010011000000100000011100011110001000010000000011010101101001101111001010111111001; 
out502 = 128'b11001001001001011101000000000001101011100110011000011100010111110101100110011001110100000001000110100011000101010110101000001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out502[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out502, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110111011001000010010011011100111101010010000010110111111100100111100001110100110110101001010110101000110110110100001110010; 
out503 = 128'b10100100001011110000001000001010101000000101100010010100101110111100110100010101001010101111100100001011000111110011010000001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out503[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out503, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011000010110000011001111000011100111111101110010101000110001110001000110011100110111101010101100100110010010110001110101111; 
out504 = 128'b01010101001111011010101010011110110011101100000110111111111010100111100100011000011101001011011001110110001010010000010111101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out504[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out504, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000000101010011101100101111101000011000001000110100001111000101010011111100101110011000100111011110001111010110111100111011; 
out505 = 128'b00001011001111001110001000111110011010110010010111110111010011110111101100010001100100100100000100101110110001111100101111110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out505[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out505, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111111100111101001001000011010000010000010011011111001100010101101010100011111010101001001010110011111100101101100101110011; 
out506 = 128'b01110111001101010001010101001100110011000001101011111011011001111110001011100111010100100110001101110010000100101100111110111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out506[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out506, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101011100011000101100010010010011001001011000001000111010011011101000001000100110000010000111001110010011100011000010100011; 
out507 = 128'b01101101101101011111111100001110000010110101100100111000010110111001100011010100011100001011001010110101100110111110011000110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out507[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out507, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001101000111010101110001111001001000000011111011001100011111001011000011001010000011011011101110000111100000110001111111101; 
out508 = 128'b00110010101111000111110101111100010111110010010101101101010010000011111110111010110000001110111000100001010010101010010110000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out508[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out508, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001011011110000101000000101010000001001100101110100101001110001011001110010010011001110101111000101110110100101000011011010; 
out509 = 128'b10011101100101100010010010110000110001001111000001011001001101001111100100011010111111101011001110010000001011000000010011001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out509[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out509, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101010100010111100001000000100011111110000100011100111011001000111111100100110111001000011000111111111010001111110011100010010; 
out510 = 128'b00110111000001000101110110010100100001111111101010010111110110000001000100100000110101100000011101001101010000100010101010100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out510[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out510, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010101001000100001110111010101111111010011101110011100001101011010111101010110000110000101010110110001000001111010110110011; 
out511 = 128'b10010000100000111101010111000011011000111110110111101110100101111011100010111101101111010100110000100111111010001001111001101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out511[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out511, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011011010100111011110010100111111010001111010000001001000000100011101100100010010010100000111000001101011001111000000111111; 
out512 = 128'b11100110110110010111101010100000011001100100010100111001111000100010110010011011110101111111110100011011001100111110010101110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out512[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out512, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000111101011001110111111000010111110001100110000111011111110111001000011011100110000100010111010111000110011110110111000110011; 
out513 = 128'b00101000011010000100110101000000010001000010011100101001010101011100110101000010001100000110011000110111101011111101111111110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out513[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out513, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010100011110110011001111000010000111011111001111010001000101111111100101111101110110101010001100110011000101011011110111111; 
out514 = 128'b00101110001110011010011000110110100001010101111000011110010001000000110001010100100101110010110110011111001010001101101011110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out514[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out514, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100100111001110001111100100001101100010101001010000100011001011000000110110011011100101010011110001111000111111010110001001; 
out515 = 128'b01000101010010111001000110100111001100000011000110100001001011000101100111110111011111110111000101111101100001000000100111100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out515[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out515, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011001100111101101101000101111100110111111011100100010101100100011001000101110000101101011001001001011101101010110000101000; 
out516 = 128'b00111000101001101101010001011111011000011001110010110101011100110100111100000001110001100101010010111001010111111011100011011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out516[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out516, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001001010011100010001000010001010010010100110010010010101000011111101110010000110110001000010001000010011111100010001111001; 
out517 = 128'b10000101000000111110100000011000111110011101111001001011100010001101110110011011100110110111110011000000110001010101001010101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out517[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out517, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010001110001010100000111001110110101010011111100111110010101111111100001100110001100111001101111000100001110000001101010001; 
out518 = 128'b10010011000101101110100000001100101110110110011000000001100011111111010010100010111010101111001011011100101111101000101001001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out518[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out518, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110101111101000010000001010110100011100100001111001001000000111110111101100010011001110010101101000001010101111110011101000; 
out519 = 128'b11101011010110000100100000101101111101000011010111011001110110110101010011010101010111101111000100001011111011011101110101010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out519[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out519, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101010000011001011011011010101000000101000110000000001001000011000010010010011011011011100111111111100000001000100000101010; 
out520 = 128'b10110110001111111000111001111010001001001110111110111111110111101101010011101101110011000111110100100111100101111100101011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out520[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out520, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011111111010110100101101100100111000110001101100000100011011101000010111110011110101000000101110000101111111100111111101000; 
out521 = 128'b01111001111111001000110100100000100100000111010001110100010101110110101100101000001000101100000010110101110001110000011011100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out521[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out521, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011101100100001111101000110011100101101100100111100111110111010000001100000100111001100001101100100110110011111110000110110111; 
out522 = 128'b11001100001101011101100000111001010101001101011001001010000011101001011000100010000001101110011000110110001011111011010001010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out522[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out522, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000101001010110001111011000110000111100100100001101010000111111000010011011010100110101101100000010111000111011100011000110100; 
out523 = 128'b01101110101110101000011011011111001101000110011100001010010000000000000011110001001011110011010000111110110010010101101000001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out523[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out523, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001111101000101100110010111111111110111011001000010000011000011000111100001110000011001010100000000000111000010110011101100; 
out524 = 128'b00001010011001001111000000011000111001100010001001010011101001100100111110010111000101111001101100110010110111001011110010000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out524[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out524, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110110000100001011111000110010111010001001010000101110001111111001011111010101010010100010111100000110000101101001001111101; 
out525 = 128'b10010100010000101110101100110001010110101001000101001100111100010010101001011101101110101001110101000001011000011011100110000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out525[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out525, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001000011101000000100100011010011100110100110111001000000000100010101011100110101001011111010001010001010101001110001011000; 
out526 = 128'b01100100001000100100111100000111100000111110100001000100100110101010011101100001111001010011000101010000110101111110110010000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out526[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out526, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110000101010111100000101110001011111011101011101100001011110011011110000110101000111001100000100111011000111010011100100101; 
out527 = 128'b11000110110010101001011011001000110010000000111010001001010110111101100101111111110010001101010011110110101111011000001010101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out527[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out527, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111010101101101110001011011001000001111101111100011001100111000000111101110110101010001101001000000001100000110110011111000; 
out528 = 128'b01101100110010111010010010000111100101100001111001001101111110000000010001100110011000101000111011111001111110110110101110100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out528[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out528, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101011101001000111110011111111100110110110100111100101111011101111001101110110110000100100110000111001011110100101111001010; 
out529 = 128'b00011100010000011001101000111101000000111111101010001001101101000000110011011000010100111000110010011110000001100001010110110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out529[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out529, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101000011011010000111010101010100101011111100110001101011110010100001100101110010001000001100010010001010100010101000000011; 
out530 = 128'b10010000100101010101110001100110111011011000110100101000000100101001110101111100111101100011110011110100101100011011011110011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out530[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out530, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011010110111110000101100101110001011101110010011100001010010001001110100001100100001010011000111110100111101000111110001101; 
out531 = 128'b00011000001001001101101111110111011111001000000110110100100101100110011111001111001011100000000010010001111010100011100111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out531[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out531, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101000010001010000100100001100010101000000101010110001100000111101001010100100010000000001001110101110001101000100011000010; 
out532 = 128'b11111101110001110011011001010011011000001100001000101000101100110101101100010111110101011111110111011000000011011001001100000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out532[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out532, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000011110011000100011101111001000000110011011010110111111110111110000111110110110011001110011100100101110100000110101100100; 
out533 = 128'b01101001111110101000111100011101001110011001110010000100100110001010110110010110111011101111111110011110010101011111110001010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out533[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out533, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100000011010101000100011111111111110111001001010001011001001001101010000011101110000010100110101010100100011010101011100101; 
out534 = 128'b10100100110111111011001100001011110110011110110011101000001110110101000010101101001001010100010101011010100111000000100101100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out534[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out534, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001100000010110011101100101100101001101001010110011111000100100010111010110101100110101101101001101101110000111000011011011; 
out535 = 128'b00011000011010000100100111000111110101101101110110001000110111111001110010110111001000011101101111010011100111100000111110101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out535[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out535, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100110100001100101011011010010000011101101010100011010000100001111100101000000110110011101000110111110101000010110100110110; 
out536 = 128'b01100001100011110000001000101111000001010010101101100000010010100011111111111001000011000010110101101111100101111110010101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out536[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out536, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101001011110111001100010100110110010101001011110101000011010100000010100111010110100101100001011001100101000000101101101000; 
out537 = 128'b00000001110110101011001011111100100100100010000101101100111111011110001101101100010110111011110000011110001001000111111110000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out537[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out537, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101110011001110010101111100111001110111000101101111001110011011000101010100100101101111110100100100001100101001010110010100; 
out538 = 128'b01011110110111101000000000110111100101011000110110110001000010001010011011110001011110101010111100110001110110111010111010011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out538[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out538, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001011000001101000010000000111100010000001010001010011001010011011011001011001001100001100010100010010011010100100001000001; 
out539 = 128'b01110101000001000111001000111001000110110101111100010010001111000001110000110101011110010111000100110110101101110010101000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out539[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out539, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000010110100111011111110000111110000000011010101000110001000001001000100001100000001000111011111000101011100001101000000010; 
out540 = 128'b00110000011110001101100010111100001110110101000100100101000011101010001111111100101011000010100100011110000010111110110000100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out540[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out540, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011110101000110010101111011001111110011111010101001000001101100001111010001101110111000101010001111110101101010111110011001; 
out541 = 128'b10011111000101011000011101000111000010101101001011101110110010101000100101010111010001010101100000101010111000110110001101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out541[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out541, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001000101001010011110111000100000010010111000010011011000000100101010111101100101011001000110110100111001010101111111010010; 
out542 = 128'b01101111011011101011011010011111010000101101111110111000110110011100010111010010110010100101000011011001100010010101011000110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out542[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out542, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101100001000101001010001011101101010111101011100001100001000000000000000111000111111011110111001000111000111000000110110000; 
out543 = 128'b01011100011101000010100101110101000000010100110110111110001000010101110011110010000110000000101001010000101001111011001111110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out543[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out543, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000010001100101011011011001001110101111010100100010110011011100000100100111111110011110100110100011010001100111101001011111011; 
out544 = 128'b10010110101100001111000111110010101101101011111101110000001001110101111101000100011000110000110101000100101011111101100100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out544[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out544, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000111000001011000100011010001011110101001011101010000001110000110000100111100011001000111101101010111010111101101101010000001; 
out545 = 128'b11000110000011010001110111101001101011011010100011111101001011001110111111000010000110001011111111010111010001110011001110000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out545[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out545, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110001101110111100011101011000101011011101010101011000001000010000011000111110101110111011101001111000001001100001101101000; 
out546 = 128'b11011101110100101010010101110000011101100101101001010000101100011011000110100000101011011110011010110011101101000101010001100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out546[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out546, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101101011000000110001101110010011000101010010111101100111000100111010101001100010101100000011100000111001010010110000110000; 
out547 = 128'b10101000110011111010110101000010110100011111111110111101110110111010001001000001100100111110011111110110010101000100001000111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out547[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out547, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001010001111101000111100000011011111011010011101010000000100101100011000100001100000100101010001100100010110111100000111011; 
out548 = 128'b10111111000010001110000000000101001011101111011100001001100111100000011110001110010011111000100001011010011000011100101111100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out548[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out548, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110011000100111101001111101101011000100100011111010011100001011110101100101100010110111101111100001001101010001010001000111001; 
out549 = 128'b10100100001001011101100110101000001111100101100110010111110010000100011101000110000110110000011010110011000000001001101000100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out549[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out549, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110000010100100101010000111101000100011110111001001011110000100100111110100100110111000011111010111010100100111010100100001110; 
out550 = 128'b11001000110111011011110010110001001011001100101110001001111011001011110101010001111111100011100100101111010001111111001110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out550[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out550, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011100110110000011110000011110000011010000001010101001010010011000111110101100000110011010001110101101000001000100001001100; 
out551 = 128'b00110001110111011000011100010101011101001100010110101111010000011000101000100001010010000101001110111010010110011110101110010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out551[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out551, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110000101001111000101110000010100110110100111101111110001000000011110010010011100111001111000000110110100010110100010011011; 
out552 = 128'b10101101101000101100110110110000110010001101010010000111000001111101011111110000111000011111011011001010001110011010011101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out552[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out552, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110001011101100101001010101010001101100101100011100110110010100011100000111010011001110101001100010110011010001100111110101; 
out553 = 128'b11010010101011010111000011011000100000011101101000101101111011110010100101111010101100010110110010110100001011001100101000111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out553[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out553, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111110000011110010100100101000101110010101000000011010111101110101110111101110111101110111001010000101110011001010001101001; 
out554 = 128'b11000010101101010011101001010000001001110011011111010010100001110000001100111101000001101110101010111101011011011110110001011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out554[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out554, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011100111001101011101000110000000001111101100111001011101001101110001111100001010011010000011110000101001111000110110110111; 
out555 = 128'b01010111110001000111010010100000101101101100110111111000100011100010000101110100101011010111100101011100011100100110111011010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out555[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out555, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101111110000001010011110110111010111000011101001010000000000101100011100000011101001110110011110101001000000010001100101000; 
out556 = 128'b10000100011100010010110010101101000111110101001011011101011000111101000110011000010101111100101100100011110101000001001111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out556[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out556, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010000100110111110111011001110000111001010111110000100100101111001000110110000110000111100001111110011011111100110010010011; 
out557 = 128'b00111001010100001110011011110011011001101001111001111111000101100010111010110110100011110111011000110110111001001000100001111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out557[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out557, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010011100000011100000000010101011000011110001010001000110100010010110101010111100010010110111111000001101110011100010111101; 
out558 = 128'b00011111111001110111001101001000110100100100000110000100101001011111111111101110010111001111111001110110000111001101000000000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out558[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out558, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001000010010010011010111100100011010111000001011111010100110011010101111110010111110100001110011010101101000011010000011110; 
out559 = 128'b01111110110101000000000100111111001101010010101110111110000010111011101100110000001111011010011011111010011110001111000110100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out559[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out559, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000101101011100010101100111101001101111101110011100001100100000000001101011111001100101100101011001100000110111010011011000; 
out560 = 128'b10010110001010000110000010000110011110100111000110111101010010101111111100101001000010101110011101000111000011111100001010101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out560[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out560, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001010101100110000011001111010110010010111010001100000011101111011001100011001011100011110101001001010100011010100010000000; 
out561 = 128'b10011010001111101001011010100110011010101101000001100100011000110011000100011001101010110110100101110011110000000111101000011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out561[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out561, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011110010100001111000110010111100010100000100001000100001100010101001010011001000110001010010001010101110101101000001110111; 
out562 = 128'b10111000011101111010000010010110001101011010000011010110101110100001000100000001111000010000001000111110111101011100011001111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out562[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out562, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101010001110101000100011101011100111010000111000001000001100000111000110010100111011011011011011011111101101001011010010000; 
out563 = 128'b00010101001111100111110101010101001000100111010111001001111100101100110011001000101000011000100110110100101011011001011111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out563[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out563, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010111011101111101010110000111111111101101000001101111110001101110100101011111100100000011000011110111100100111000101010001; 
out564 = 128'b00111111000011110111100001110110111000001011010010110111101000101101111011111011010001100011011100000001001110010110010100000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out564[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out564, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010001111100011011010100111101100010101111010001001101001100011000110101101010010010111010010010000100011110010110011111101; 
out565 = 128'b10101111000010110110100110000100000010010011101000010000000100100111011010010001111110000011100111100100000011010111111010011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out565[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out565, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110101100001010001010011110101011110001101010001001111010100001101011001101000000000001101100000010001100110111111011011000; 
out566 = 128'b11110101011000010101000011001000001100000101101011001011000111000001100000110001101111010010101101011001100001111101001100011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out566[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out566, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001010111011101011110100000010000011111010100111101100001011110000101100100100100101000001011101101110010110111101101100100; 
out567 = 128'b00110111001111001110011110101101101111010111000101111001001110111101011111110110111010101101010000001111100001010001010010001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out567[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out567, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000010100011100110110001111000100100000000100000110101111011001110111000111101011001010011111001111111000100010011110000101; 
out568 = 128'b01010001010001011000110100101101000101011110011110010101111110101110000111000110111010101101110100000110100100110000100001111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out568[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out568, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000011001111000001010001110100000111111111100011010111011101001111011011101100100010001110001100110100010001010000101101110; 
out569 = 128'b10010011000110111011001101010001111100000001000101000100001010001010110000101101001000101011000111000100100011101001110000100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out569[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out569, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011111011000011100111110000111000001111100101101010100011101111000100000101010010110000110000000011001100001000110101011111; 
out570 = 128'b00101111010001111000010001110111001110011001110011000101101110010000101101110110101011100000101010100001010110010011111000000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out570[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out570, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000101110010111001111001010100010101011011011011011110000000010101000101110011000110010011001001000111001100011100000110110; 
out571 = 128'b01001111000001000111010110001101010010010000000100101101111101010111101010010100011110001000010011111101010001111011010000101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out571[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out571, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010110010001001100111001001100010011011111001111001000000111101111100100000011101110110111010001000100000000010000100001100; 
out572 = 128'b11100101110011000100110010100100101110001111110000100111001000111011011010000111010010111000011100100100111110001011110111000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out572[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out572, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100010001010000111110010011000100110000100100010111101001010011000110100101001000000000001110011111011011011101001101011001111; 
out573 = 128'b00100011111010100011110011100100111011010111100000000011110011000010100010100111101100110011101110011100111010000111101011010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out573[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out573, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110100001110000011000100101101010100100100100111111101000110111011011110101001011011011110110010000111110101101010100011110; 
out574 = 128'b00111010000011000000001011100101111010010100101011110000001111100011100111001010100001010001111010100000000100110101111001110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out574[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out574, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011011010100110001001110100001100001010100101010111111101011000001111111111100100000100011001110010000011111010000110010111; 
out575 = 128'b11110001110101111011010001011111110111000110100111111010110101101000111000110111010110001011111011111001001110111000010011101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out575[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out575, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001010110000010111100011011001100010101101101110010011011110110001101011110111010010011011000011011000111111000010100011110; 
out576 = 128'b10001010000101101001000111011011000111101100100001110110100101001111001111100111111101101010000100101011010011111010010110000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out576[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out576, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100100101111001000010101010000011010011000011101000101100011000101010111000100010000011111000111010110010000001011110110001; 
out577 = 128'b10111000101010111011111110100010001000000011100000010100000101111101010000100111001010001011101000100011000100110101000100110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out577[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out577, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101010011010100010000100001001010101000011000110100001010101000010110111111001101010101000011010010000100111011100001000010; 
out578 = 128'b11100011011111011111111110011001111011111010000010000101010010100010011110011001111110100110000101100110010111000100111010100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out578[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out578, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000011100101101111100110000001011010100111011001100111101101000100110001110101000011001111011110110011010110000100101001101; 
out579 = 128'b11100100101010101000001110110011110010010010001000101101100011010100000011110010010000011001001000000011011010001100101101110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out579[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out579, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101101100100001010001011001001011001111000011100101111011000110101101101110111000000000110011010011110111011110110110001110; 
out580 = 128'b10000100110111100001101110000001101011110001011110100100111011111000000110110010111001110110110010010110011001111001001111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out580[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out580, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101111011010100100001011001110100010110110000010111001100110000011100000011011100000110110101011110101001001000111100111100; 
out581 = 128'b11110111011001100001101011111010000101100101000000111100000111001111010001110011011100010000101100001011010000111101111101100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out581[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out581, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010000100100110001111001011011110001011001000010000010010000110001100100011110000010111100000111010011110001011010001001100; 
out582 = 128'b00100011010100110000111100000011110100110000001010101010101101011000101101111001010000101110010111010011111101100010110101000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out582[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out582, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010111101010011111110010111010000100010010111110000110000010011110001011110001011000010111111110011010011010001001101001111; 
out583 = 128'b10010100011011000100111111001010000111000101101010110101010100100000011010111100000001010111001111101001100001011110010100101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out583[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out583, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111111000110110000100000011110000000101100000000010111010100000100100001111101000000100011010101010001011101101111001011000; 
out584 = 128'b00011110101111001000100000010000010110010101101110000001110110001100100011111101000100110100101101011111001001010000100100111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out584[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out584, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101000101111101111100000110010110011110001000010000111110010000111000111000101010001100101001001000000000111011110111111010; 
out585 = 128'b11010011011101000000001000010100100011000110011111010101110010001101010100101011010100100011111000100110101100000110010010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out585[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out585, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000100000101101000100000001000010001000000111001101011010110110101001001011101111110100111101101101011111101110010100111011; 
out586 = 128'b10111000010111111111100010010111100011100011010110000100110110011101100110110000111110001010110010000110001000001100000110101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out586[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out586, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001100000110001000001010111101011001111100001000010010100010001011110101001101101000011111101101100010111111000010011001001; 
out587 = 128'b00000110010011101100101100000000000111011001101110100010110000110000111000000110101000000100001101000111010110011000101101101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out587[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out587, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010001000010111100100111010110001001100001101001101011110011101100100111110001111001001011001100000110001101011110100001101; 
out588 = 128'b00111111010110100110011000110010010011000100101001110111001001101110010110111001011000001010101010111110110100010101110111000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out588[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out588, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001010001000100101111111101000110011110110001110000100101010100001111001100011000110011110001000110001111010001101111100110; 
out589 = 128'b10011100011011111111011011111101011110110110110000100101011011011010101011111100000111111000110100000000010010010011000100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out589[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out589, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000110110010000000100101101101111100111110100011011000110011110011001101010011001000111000010101010010001111100100111001110; 
out590 = 128'b11110101010110111001110001010111110010110011000110101010000010110100110110000001101001101110001011001011010110000000100100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out590[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out590, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000011100011110010111000010011011111011001001001111000111011011010110011000100001110110111000100111011001010110110000100000; 
out591 = 128'b11110001001001101100100011001111100000011001110111100011111101110101001000000100111011101111101001100001001000110001110001000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out591[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out591, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001011100111111100110111011111000001101110001000100010010100010100001101101110111101100010010000100010100111011000110010000; 
out592 = 128'b10011110101010110111100101100011110001101001110010011010110110100010101010000100110101000100101001011011010001100111111100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out592[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out592, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000100011000001100000011101111111001111001001101010000100100101110001010100101100111101010000000100001100101100001010010011; 
out593 = 128'b10101101110101001000011101010001101000101101110110001001011111100010010111100111110010110010100000010100111110101011100011110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out593[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out593, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000000110001010100100111010011101010011111100011111011101000111111100101100100110010100100001000110111101000100010111100111; 
out594 = 128'b10011101000000000001111000101001100110101001000010101001101101001001000100010010101101111011110111101101010111000101010000010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out594[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out594, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000101110101010011101010110101000111010001111111000101001000000110010110100101101101101011100111111101101110111011001111010; 
out595 = 128'b10011100110010011100010100000011111101101001101100110011000001011110100111000011010000001100100110010001010111001101111101001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out595[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out595, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111101111010000000111100111100010100001110111001100100010000000101001011011010111000001100110100011110010101010100111101100; 
out596 = 128'b11000000000110010011110001101100000111000010110110111100000010101111110000010001000100000010011110000001100101010101111010010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out596[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out596, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010011000001101110000001001110000011101110100001110101011010001000110101010011110111110001011001010011001111100110011001111; 
out597 = 128'b10100000101111011100101111100100011110101100000000110001101100000100011111100001011000001011111001110111011001100111101110110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out597[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out597, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010001001000011101011101001011011010100001010010101110110111010011000000110110101001001110001011011000001110110010110011111; 
out598 = 128'b10010010111100111010000101010111100111000111011001110110000001101101110010111001110111011100110111100001001100001111100010110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out598[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out598, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111011100110000111010000000001001011010110110100110110010010110011001010100111010100000110010101001001010111010100101110100; 
out599 = 128'b11011001101110101100101001010001110100001100110001011101001111010010001100011101001111100000011101011001111110010011001111111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out599[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out599, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011001100100110111110010111100011001101001011011101101000111101011001001001001010110010100010011111101111100010111101110001; 
out600 = 128'b01110001100110011000110100011010000000011010011010100010101110011011000011101010111001010000010000101000100111010010111011110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out600[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out600, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100111010111001111100110101110011101100001011110001101111101001101110011110001011011000010010110100111110110000100001110010; 
out601 = 128'b10100001010001111101011110001100101011000010101000001001111011101111001101101100011011010110110010100111010111011000100011100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out601[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out601, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000011010001100100100111011000011000001101101111010111000100000000000010110110010110010010010000111101011000000011001110101; 
out602 = 128'b00001111010100110110011011010000001001100000001111011011001110111100100101100111001001101100111011001100111100110000111111011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out602[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out602, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100010101011011011111010010101011100001101001010101110011000011111000110011011000101111010101100111010010110100111011101001; 
out603 = 128'b01000110000000001010110001111101110100100001100000010110010000101001011001100001100001111001001101001100111100111011101110110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out603[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out603, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110110110011101101010001001001110010001101011011101010011010111011100001000100010110000101000010001000001000111110001011001; 
out604 = 128'b01001010110101111011010111101000000000110010000111100001111101010110010000111100011001110110100011101001011000101000000110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out604[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out604, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111011100111111001101010001010111101000101101000011101110001110101000101010000000011011111010101101001001100100111011100100; 
out605 = 128'b00011110110010101110010011101000000011000111000000001100100001001011111101010101111000110110011101101010101001110000111111110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out605[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out605, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001011111000111011011110011001111100010000100110100110010001101000010001101111000111000010111100100010111111100111100111011; 
out606 = 128'b00100010000110111100101100100001110000001111111111011110111011000001101010110010001001110011100100011001001110100100001101010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out606[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out606, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011100011100000010110001011101100000101111000101110010110111001011101011111011111010010001011110110010101011101111000100101; 
out607 = 128'b00000101100101011011000111100011100001111100101110110001001111110001101100110101001101100011000100100010111110010110100010001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out607[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out607, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000001100000011000011100000101000001110111100010111011001000010111100111101000111011001110011111010010000100110001101111001; 
out608 = 128'b11001101001101111011010111111110100111101110101111111010000101000110000010011111110101110011011001110111101011101111001111101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out608[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out608, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111100001001101000101010100110010000101011100000111101000111111010010011011011100001100110111001101001011000000001011101001; 
out609 = 128'b01001110000000000001110110011011000111001010111110111100111101011010001000110111001011011001000011111010110100010011000010001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out609[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out609, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001111111010111100001110100110100011010000110000011001001110110101001110100000001101000111000110000101001110101101110110101101; 
out610 = 128'b00111000010110011000001110001011000110000000011000110101010100000011011111110101011100110010101010100010111111110110000100111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out610[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out610, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000000100001001011111101001101001111111001100110101010010011011000010010000110010000010110011010010101100111111011010101010000; 
out611 = 128'b11000110000001100100101111100110011100111001010111100000101100101101101101000001010000010111001101101100111000101001011101110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out611[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out611, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101000010000000010100101010001011111001110010000101001000101000010001010110100100001111101100011101100111100010001111101000; 
out612 = 128'b00010111101111101110101100001000001101110011100010001011111000011101110010111100110010111011010111100011010000001000110110101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out612[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out612, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100100011100111011100111110010110010101110011110111000011100101011100011001010011111011101011000011011011101101001100110110; 
out613 = 128'b10010100011000111111100101000011000011001001110100100011110010011101100111101110000001000111100110001000000000001110111111010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out613[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out613, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100000100100001011000111010011100101011111110110010101010000101111010000010010110100010001111100010110110001011010011101101; 
out614 = 128'b11000000011111111111010000100011001101001100100010110101011010000010100101101110111011100100001000001110000001011011101000110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out614[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out614, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011110011001101101000010111011100000100011001101000001000111100010101001110111010101110000101101101101011100000100000101001; 
out615 = 128'b01110000110111001111000010110101100010110000101100011110100111110011100011110111110100100001100110101101111010001001110000101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out615[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out615, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011011010011100011101000011001001001000111011100101010001010110011111011001111011110001011010011000111100000000110110111100; 
out616 = 128'b00100111011010000111100011000011110011011011011110111011111010100111100001101111001001100000000101011101010100110011101010100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out616[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out616, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010110000001011000000110001011011111101001011101100011100101001100011001101010101111110111110010101111100001110100010111111; 
out617 = 128'b01001000001000110100001100010000101010001100001000001101001101011011100101100110111011100010000110101011011011011101100111000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out617[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out617, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100101011000100100101100111000101011100111000001101001011110111111100101001100000001001110101110000100001010101000101110000; 
out618 = 128'b01101110010011010101111100110011001010010110001011110100010001000110111011010100110011010101101101100010001111001100001010011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out618[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out618, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001011001101111001001001100011101100101110001000011110101001111001010111010100000011111110001001100110101011110111100011001; 
out619 = 128'b01000101101010001011111100100110001100101111111101010100100110111111011110010000111000101100001010111011101000001110100000010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out619[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out619, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010110101111000001110100001110101010001101011101001001101110001010000110111001111101011010010011110110010111100000111011100; 
out620 = 128'b00101000110111001011000000110001100011111101101111110000111011100011000000000011011011001001010000010100010100101010010000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out620[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out620, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000100011011000101100011000001001011000100001101110000011011101101111010011111101101001011011000100100000111111110011001011; 
out621 = 128'b11011111010001000001101011101101101000000000100111011000011000001110101111011111011010111001001001101111000100110001111000111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out621[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out621, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100101100111000011001011110110101000101010101110001101011011010000000110110100011111111010010100010011100010110110011010111; 
out622 = 128'b11000010101000100011010100000011000011000010010101100000000101001100110111001010010100001010111110001101011111011111111101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out622[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out622, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111111111000100000001001011001011001010000000101100011011000101111011111101011011010010000111011011101100110110111001111000; 
out623 = 128'b11101010111000100001011000010001101010110110100010000001010010110001110111000110001000101110100100100100001111000111111110110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out623[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out623, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000111010101011011010001000101001010100100011010110100001001011000001110011000111000000011000000001100011011011011100000110011; 
out624 = 128'b11001011111010000100010001100110101011100011011001110101100101010100101110111110101011110101110110011011101010010010001100001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out624[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out624, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001011101100100001111011100010000101111111001100000100110101001000011011000110000001111011111000011001001000001110111111001; 
out625 = 128'b10001000011001001000111000010110000111000000101100011011011001101111001000110101000011001010101010110001100000110100011001011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out625[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out625, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010111100101010000010100000001100010000100000010110111111001011100011011001001111100110110010010000111111100100110001110110; 
out626 = 128'b00100000110110111101110010001000110101110000000101010011101110001110011110001100010001111011000110111100011000010111100011101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out626[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out626, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001011000111011010100100000001101100011111110010010111111111010001000110110010011101111010101010011111100011001111111001011; 
out627 = 128'b11101101110110000000011000011010011110100100001110110101011111110001100100011001100100101100001000000100110101011101110000010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out627[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out627, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011100001101110110011011001010110011000000011011111111100011001111110111000101010000010000001101110110100100110100001001000; 
out628 = 128'b11101110110010001011101011100100101010111111001110110011010110000100110000000001011011000011111000010010101101111100000111011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out628[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out628, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100001111011010010000111101111111110101111100110111010101100100011000111010010010000000101101100001100001101100100011011010000; 
out629 = 128'b00100110010010001000010000001010001111101111001100011100000100001101100110100000000000000010010010001110110001100110010001010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out629[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out629, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001001111101001101100001001000100110010001110010101000010001101000000100100110010000001100111001000011110110101000101101100; 
out630 = 128'b00000010010011010011010011011011011001100110010100100111100001100100000011010111100111011100010101110000000101110100100000110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out630[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out630, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100010011100110110000100110100101101111101000111110010000001000111111101111100000100001001101110010010110100001100001100100; 
out631 = 128'b10101100001000110000110110110010110010000110111110100110101100011100000101101011110100001101101110000110110110010111011010001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out631[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out631, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101011010011111011101010101010011110011011111000101010011011000010111000101010000000111101000101111010001110001001011111101; 
out632 = 128'b10011000110110000100000010100101101010001001010100101111010010011001011100000001001000100011011110110100111001100100000001001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out632[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out632, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110111111010110101010000001011010000000001001011100110101110100111010001011100011111100011001011111110111111011101111110010; 
out633 = 128'b01101101110000100010101000101011100010111010001010001001111110100111010111001111000010001001100000001010100011111110101110101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out633[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out633, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000100110000001111101111111010100110000110100111011111101000000111000001000011011011011110010100111001000101100101010010110110; 
out634 = 128'b01001110111010101111011110001010101100001101101000011001100101000111010101110111001001111011000111010100101011110000010101010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out634[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out634, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000010001000110001111111110000001101100011010000011101100000111100111011010011000011001001101100110110100110101111110000100; 
out635 = 128'b01011010111110111010101010001111000101101011000011101100001011111100110100111011101001111100000011101101010000000111110011110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out635[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out635, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101011101010111010110010101100101001100000001000101000010000000001100110000111000111000011111000111010111110011010000100000; 
out636 = 128'b11001111000110000010000001011000101010001010110100001100111000000101111010010001000111001010100111101111111101011110110100100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out636[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out636, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100100110001100000101101010000111010100110000010011010000001010101010000100010010011010110001000011011101110010101001101001; 
out637 = 128'b00100010100101000100100100011110111001101101101100010000111001100100100111010101110001111001010010110111001100011000100101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out637[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out637, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001000101001111101000001110001110111000011000111100111100010100100110101110111101010010000011011110011010010100100011100010; 
out638 = 128'b10101100111100011010001001111111101000001100100101110110000000001011101111011100000110110011101011111001110001010111111100000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out638[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out638, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001110100111111001100000001100100011011111011110001010001000001100010001100001100100001111100011010001011011100110101110011; 
out639 = 128'b01011010100101001100110000001111011001010000011100010111011000101010011100110110110010111101011100110110110000001101011111110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out639[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out639, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101111000110111000100000011010001100010000011110011110111100101101010001110010000011111011111000100100111101111010101111000; 
out640 = 128'b01011100001110011110001011101101100001100000110100010001101000000101100101011000100110111111001100110010000001001011100110100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out640[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out640, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000010111101101111000101011110010111111101000010010010010001100101011111110001101011110010101101010011010010010101110101110; 
out641 = 128'b11101110100100001111000111110000110101101101000110000110100101101110100111111001110011100000001000110111101010101110110001100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out641[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out641, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100001001011000000110100101101101001001001010100100100011011110010101101010011011011011110101110101100000111001000100000110; 
out642 = 128'b00110110100000111111110001111010010100001010110111010010100111000001000011111001011001001100001100000111111011111011010001010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out642[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out642, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001011010110100010100111000110101000010010110001010011001101001111101100011001111110000110101100101101110101001001101011000; 
out643 = 128'b11011101110100010111010101000111011010101000000000011011100001100001101000010110111011111010001101110000110101101001101101000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out643[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out643, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111011111010000011000001011010011000110110011001111100000010111011111100100110011010000100101101100000011000111111011000101; 
out644 = 128'b00000001010000001100111000000101100000011000100101010001001101011000001101100000111000100101110010001001101001001110101010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out644[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out644, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101000101101000101100100010000000110110111100110000101011101010100110111010001111001000101111001011110100001011111101111111; 
out645 = 128'b00110111001111010011110000001011000111011111110001011010010001110001110101001110000010110000110110001000110001001111010011100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out645[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out645, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100001100100101000010011011101000110010110000110010010010010000110010110100101101111110101000110100100010011000101000001111; 
out646 = 128'b10010011100101101101000010110100001101011101001010010110001101000111001011111001011000011001101011011111000110010000001000001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out646[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out646, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101100101111001010110101100010001101000010100110010001101110010101010010001100000010011010000010110100101101011110001110111; 
out647 = 128'b00011011101001000001010010011011101010000011000100011011101100110000000011110000100000010011000110000001111110111011110110001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out647[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out647, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011111111000100000110011101011110000011000110010100000010001001100001001001011111001100111111011000110000110110100110010101; 
out648 = 128'b00010011001101010011000010101101100111110010000010011111010000010100110010010101001111000110110001101101000110110000111001010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out648[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out648, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100000000011011111110011010001110100101000111100111011010001100101110000010011101101111000000100000001010000111000001000011; 
out649 = 128'b10100001001000100000101111100101111011000000001110000000010111011010001001111111110010011100001000110001011100011001001000011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out649[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out649, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001101110110010111011011110110001101001111010111000110101001100111111001101101110100101110010000001101111100010000000111100; 
out650 = 128'b00111100001011011011111001110000100111010110110101000010001101011101001110001111001110011100110010101100010111101110111101101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out650[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out650, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001010111111111000101000100001101110101101001010100110101000111000000001100000111110001001011001110010000101000000001100011; 
out651 = 128'b00010011010111100010010001110010001011110011000101010101000000111100010001001100101110101110001001011000010110010110000011110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out651[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out651, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100011100010000001110001000011111110011001010010100001010110111100101101000101000011111011100000100001001000010000101100010; 
out652 = 128'b00100101100101100101111111010110000001001001010100001010101000100001001010101110110011110110001111010000011100100110010010011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out652[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out652, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100101110010011000011111100111101111011100110010101111111111101100101100000000101111011111000011000110000111000010011011001; 
out653 = 128'b00100010111110001011110100010110001100111011100111011000011010111011000010110000010100010001100110001011010101101111011011100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out653[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out653, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000000111111100100000000011011100000111101011011110011101111000010000001011010100001000100010010100000001000010110110000011; 
out654 = 128'b00110000111001010100000001101000110010010100111000000000010010110101111110010110110101100011010001101100011010010110110000111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out654[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out654, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101000111111100001000011101011100100001100110011000000110100001011011000001011001100111001000011011011110011110010011001110; 
out655 = 128'b01011010011001111010111001010010100010011010000110010111000111001000000010011010110111000011010100001011010010110101011100000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out655[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out655, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100010111111101110010000011001011100001101010100110000000111001001001101100110010011110101000101011000111010110101000001111; 
out656 = 128'b01110011011100111000101011100110101011110110010010000010101000101110100001110100010110010011000011101001100100100010000010101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out656[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out656, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011100111100001000111110100111100011001000110101111110100000010101111001110110011001010011110001010011011001000011000110011; 
out657 = 128'b01001110000001110101101110100110010111111101010110001001010010111101110110101000001011000010010111010010101110100000101100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out657[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out657, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110100110011011111111011000000110001000011011001111001111101010110011111000110110001100100111001011111111111000001010000101; 
out658 = 128'b00110010100000110101110000111001101111100010001110010101000000100001101010001111010000000000110000000001000100011001010100011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out658[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out658, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010011100011110010101010001111101100001100101101001101001010011110111000010100001000100011101000100111000010001111111011100; 
out659 = 128'b01010010100101100010111001001010110101110110111000100000011011100110111000100101001011111100101100010010010100100000001100101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out659[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out659, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100011001001110011111000101101000101101110010001101101101011011101111110101011101100010101011010101010110011011000000110111; 
out660 = 128'b11000111101001011000110000101001001100000100111110011010010110110010110001110101011010011101110100111100110000101111110010111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out660[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out660, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100101010100111101110111000011101010001000110011101111001000000011000111010101100111111111111000100000000000011100011110010; 
out661 = 128'b01100000000010101010010101010011010010010110001100100100100011111100010100011000001010001001001111001010100100111010011000000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out661[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out661, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011111010110011001010111111010111101001101101010011011010100000000101000001010101110000000001010010101100000010101011101001; 
out662 = 128'b00100100000011100101111100010001011110010000010110101111010100001100010010100111110110001000110100011110101101100000001011111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out662[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out662, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100100101111100011011101000010100001001010101010110000010110000010000010101000110011111111000010110001000110001101001000100; 
out663 = 128'b10111110010111101011010001010011001111111110100011111101101100101000100001000000100111110001001000111111110111110101110011110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out663[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out663, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100010010010110000101010010000010111101101001001001000011100101001001011000100001100101001000001011110100011100000100111011; 
out664 = 128'b11101011100111001101001000001100010101000010111100011110010010010011011010011100101001111011010111111100001110010100101100000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out664[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out664, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000110010000000000011101101001011101000011100010111000011111011010111110010101100101001001001011001110101101110000100111000; 
out665 = 128'b00011111100011111101110111000010100111011011101000010000110000001100101111110100101100010001001011011101101100011000100001100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out665[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out665, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001010101001100010001100001000111010011110100110111100001010000000101000011101111010011001100110011100010000000101001001100; 
out666 = 128'b00000000001101001100100011101010101101101101100001101001001100000010110101000011001110000010011010000000000100111101110000010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out666[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out666, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001001100111001101001010100011011110111100111100101110010000010110011111100011011011111111010100000011110011001100111110101; 
out667 = 128'b00011000111111011101000001010100100000100011111000110111100101100111010110111010101010100010011011000001100010001010110010010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out667[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out667, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000011000011100001010100000001110011110110110101000010010000100001100110010100001010001000011101110010110000001011011100111; 
out668 = 128'b00000010011010000101101011001000101000010101101011011001110101011111100011001101010101111101000110101011101111101100001011001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out668[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out668, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010101011101001110010011001010111110111111100110111111111000010110001110001010111111011011010010110001111110011010000000111; 
out669 = 128'b11110001110011100010010110111000111010001100001101010011001100110101001001111000011011001011111000010101010000011011111111001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out669[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out669, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010000000100101101010010000110000010110100110001101111101000001000010111100111100100101010010100011100011101011000100010110; 
out670 = 128'b01000101010101100110110101100001010011101001001000010101110110110100000000001110011000000100001111100110011110001000011011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out670[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out670, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001111100100110101000010010011100000001001010010001010101110000100011111111110011011111100010000010000011100101110010101101; 
out671 = 128'b10101011000001100100111010001001010110111111001011011000011001001010001110100011001100111001011100111100110011001100100011001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out671[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out671, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110010011011000101010111010101100011110111100100110001101001101011000001111001001010101010000010011011000100111111111111111; 
out672 = 128'b11000110011101110010010110111000010110110001001001101111101111000001010100011110011010100000010000000101100111111001000001110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out672[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out672, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001100100111111110111000001111011111001000110111111011111010100010010110001101110110110100100110011100011010010000100101110; 
out673 = 128'b11101101001000110111111100101000001100111011000101000000001101011000111101011100010111111100011001100000010001110110011110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out673[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out673, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100000000110000101000110101100011111001000110011001010000000110101001110111101000111001111111100101011011001101010011101000; 
out674 = 128'b01010110011101111001101010111001101110110111100111111011001001111011110100101010010000110110110000111111001001010011110011101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out674[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out674, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011100110111101010101000010111010111101111101011001111010101000101100100101001111100110010011001101100110001011011010001011; 
out675 = 128'b00101010101111101001100101101010000110000111111001000001010000011101000110000010011100001100100101001001011001100101010100111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out675[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out675, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001110010110001100101000011100001000011101000011111001110000001111000110100100000000001100100011001100101000100000110101010; 
out676 = 128'b00010111010001100000010100100011110111111010101001100101001001101011001101001010001000100111010001011101100101011001000110010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out676[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out676, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011011001010010011110111010100110110000011011110111110101110100111100001000110001000001110111100001111111111001110011010101; 
out677 = 128'b11000101111000110011111001010010000111111100000001011000110000011100010011110110101101010000101010011101111100110100110101101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out677[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out677, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010010111011100001011111011101001101000110001000011101010100101011110100110001111111111110000010000110100110011010011010010; 
out678 = 128'b01110010101000001011111000101101100100111010101001111111101101000110001001101100011101100000011110101110000001100101111010000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out678[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out678, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010111100000101100011001011000000010001110000111010101100100001011100000100001111111101110111010000010100001110110000101110; 
out679 = 128'b00100011111111101100100011001010011111110101011110000011110001010100011010000101111011110110100010010101101111100111001100110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out679[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out679, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110010001011000001111000001010101011100000011111010111110100000100111100100001001110000111001000001001000101101101100110001; 
out680 = 128'b00011110001111001100110100110000100011001100010100010100101011101101000110011110010011011111010101000010000110100111011011010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out680[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out680, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000110011111111001011111100001100100101110000000011011101101111100110010000100000101001101111110010001101001000101010010100; 
out681 = 128'b10011110011010010111110011000010100011101001111000111011110000001011001010110101001111110011111010111010111111111110100111011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out681[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out681, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011111100001101111101100101110111010101100111110101100111001110111000100000010010101001011111001001100111001101101011001001; 
out682 = 128'b10010011001001000100010110010100000101100001101000110111001111100010010111001001111110101100001111110100110111101101010010100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out682[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out682, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001101101111110010100000111111001100000110010011100011101110111100000101001111011000100010011000010011110111011011100011011; 
out683 = 128'b10100010011010010111010101011001110101100100101101001110111100001110100010010100111101100000000001101100101001101111011100010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out683[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out683, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001110100100010101111110100111110100000101101100001101101101110011001000001100101010011100010000010000110011000000001110101; 
out684 = 128'b00100010010010010100100101101001101010011111110010111100101111000000000110001010101100001110101110100101110010100111000111011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out684[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out684, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101110010110010000110110110111011101101111111101100101000111011011010100100111001001011000100111001100100110010111001101010; 
out685 = 128'b10110101111001100000101001100000011010111111010110010001101110111101010110100000111000101000100000110100010111111001011111100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out685[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out685, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011101101010110100001100110010010000111101100010101111010000011101010011110110000111110100100111111100001101111010111111010000; 
out686 = 128'b10000010000010110010011011100100010001001011011100110100101000111111100101110100001111110101001010100110101111000000000011001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out686[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out686, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101011110001111101000110000011101000110111000001000010111111000010100011110010000011101001011000010011100111011110011000110; 
out687 = 128'b11101010110100111010001011011100100111100000111000101010101111011010001110110000011100000100111111110001010000100001100100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out687[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out687, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010010010101000110101111110111101110100110100110001000000111010000010010001101100101110001110010001101110000001001010000001; 
out688 = 128'b00111100010001000001101010000001110010011111011000000111011001110000100110101110001110100100110000001100101000110000011110011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out688[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out688, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000111000000100010000111110100101010111111010110011110101000001010111100001000110100101000111101001111000000001100011010001; 
out689 = 128'b00001100011011000111011100100010001111100000001101001101101000000110011111011011101011000011001000100010011010000000000000100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out689[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out689, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011010101111010000110101001101010000111010111001100011101001110101011110110010010111110100100110110001110010110011110000011; 
out690 = 128'b00011101011110010010101011100110111011000011011000110011011001101111011110011001110001011001101101100010101100011010110000110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out690[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out690, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011100101101111010100100011001010001100010101010111001100001001111111010111000011101101100110001110010000000101000011010110; 
out691 = 128'b11100110001010101111001011111011100001010000111101101011110110000100010011100001011010110101010101101000001000010101100001111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out691[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out691, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001111100001111011011111000110010101110000010000001101011000001010010101100000011000110010011011001001011101001110111100111; 
out692 = 128'b11001110100010011000010111111011111111101100000001001111111100001100001000010111010000011000111111000001011110011111001101111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out692[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out692, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111001010010111100000101001110100010111101100011110000001101101010011001000101000010011100000100101110101111011101111101010; 
out693 = 128'b11011110100010111001011010001001111011101001101001110111011110100111110010101100001101100100111101010101110011100101001100101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out693[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out693, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010111001100000100001110010101000000010101101001010010101001110111101011000001111110100000111001000101101011001001001011000; 
out694 = 128'b10111111001101100010110011001010100000110111111010101010111010001110010001000010101111011100011001011011010011000001000110100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out694[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out694, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100111011000001101000001011001010011111010000100010010011101001001010011110001011110001010001110100001110100011101000001010; 
out695 = 128'b00001111010101111111001010111101011001000001011000111001010101001010101000110011000110100000011100111011011100110100101110011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out695[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out695, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110101111101011101110101011101111101111001000000011011000111100001011110101111110010111100000110011011010100001101110000010; 
out696 = 128'b01010011001101010110100100100001111110001100001001010101000000001001001111111100100000000000000111011101100010111110111100101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out696[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out696, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011111010100000011110111101110011010110111111110110011100011111010001100010000001101100000110010011001001011100100010101011; 
out697 = 128'b00011111001010001100101010001000101110110110000010100011000111110101111001111101010110110100010011010000000000101110010101010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out697[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out697, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100100010000011110110110111101101011101111110110001000001000000011000011100011011101100100111011100011001001010000010000100; 
out698 = 128'b00001100100010001110001011111000111100000000100100110100001010011001110001010011011111110100001100101101011111011011001000111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out698[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out698, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111010011011110111011100011011010001000101110111100100000110111100111100010001110010001100000110110100111111000111110101100; 
out699 = 128'b10000111111001011101011100011101010011110101001001101011011111011101010011000101110000010101101100001011011000000110111011011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out699[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out699, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111111010110001001111011111010111010010111101010001010001001111001110101000101110100010111100110000110000000001000101100010; 
out700 = 128'b01011100010110010010001110001001101110001001011000100001001110100000100011000011011100011001011000111011001111000001101010010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out700[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out700, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000110000110001100110011011000101011101011100100011110110100011010101000010101111011101111001111010110010010010111011111000; 
out701 = 128'b10101110010001101001001011001000011111100010100011101100001101000010010010011010100100111010110010000100011001010001110011001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out701[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out701, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101000010001001001101110001001100110010101001011011100101100110000001001101001001011000011110000001000101110001010111011000; 
out702 = 128'b11010110010000001011101010001010010010011000100000101001000110000100111010010001001000011110001010111101000000110100101101010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out702[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out702, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001010100101111000000001000110011010110111101100100110101000100100011101101000001100111000010010110001101011010000001110001010; 
out703 = 128'b10011010110110111010110111101111010001100100000111100100111101110101000111000011100110111111011100110010100011000110011010111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out703[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out703, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001000110101000101001111111111010011100110110100110001010100001001110010101011100000011100001000011100001101010100111100101; 
out704 = 128'b11010010010111010010000010011011101110110000101111100101011110110010101100000111011011000111001000001001110110001001100100001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out704[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out704, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000010011100001001010001010001001001000011011111000110100110111000010100101011110010000011101110111100000010011110010011000; 
out705 = 128'b11011111010000111000000100011011100101100110100001100001001101001010011111011011000000100010110101000110110001110111111101011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out705[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out705, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110000010010010011101001010101110100000011010001011100011111111001010010110001100011110100010001101001011100110010000010011011; 
out706 = 128'b10001100101101000001010101011000101011110110011000100000010010011101010111111000010110010010100110100001101100111000001001000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out706[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out706, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101111110000111111011110011111111000111011000010000111010000000010101011000001010001101010001011001110010010000100010111011; 
out707 = 128'b11010100111110011100001000000001010000100000100110111111011000110100010110100100111111111001011110010101010010101100011101001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out707[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out707, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111101111011101110100011111100110101100011101011111011110100111110001100011001100001110010111010100001011000110100000010001; 
out708 = 128'b01101111111000101101110101110001101100011110110001011100010110101100011111110101110011110100101100010111100100111001100101000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out708[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out708, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001100001010101010101110011011000011010001010011011001010000111110001000100011000111111101110001010111000111010011010000001; 
out709 = 128'b10001001010100100000111101101010110010100011100100111100001001000101100010001110101111001110101110010100110001000011111111011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out709[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out709, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010101100111111100011110100010011111101011011001001011001110011110011010111011001101101101110000011111100110000011100000101; 
out710 = 128'b10010001000001011100000010010101011011010000010101101101001100100000110010111010000111101011111111100000110000000110011111010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out710[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out710, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100010010000111110010110101101010001001010100000010101010100000010011010101111011110111101001001001101101010000001000000111; 
out711 = 128'b01101011111011100011010000001001011111100110100100000101000111111101110011011110000011010101111110101011101111110011011010000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out711[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out711, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101111001110101001010111011010000011010110010010011101001011010001111110011100001010010110110001101001000100011100100111001; 
out712 = 128'b11001111000010001001011011110000000110001000001100001000101110001010001011110000011101110110100000010101101111011011111001010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out712[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out712, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101001010011011110011011110111110011111111111111110001111001110011110011001111101110100100110001101010000101000000110100000; 
out713 = 128'b11110011110111011101111001100001000100101111011001100011011011010101101100101100100110011111101101110110010110001101101010010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out713[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out713, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011000010100111100001000100111001001010111001101111100011010111011010000011100110000111010010001111110100010011001010001001; 
out714 = 128'b00101000001001111000010111101110100011010111001011011001100101110110000000011100100110000011000100010000010110111010111010010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out714[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out714, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011001110010011001100110000111001101011100001011100100010100110001011100010001101110010001110111101010111011011111101010100011; 
out715 = 128'b10011110101011100100111110010000100001011010001001110010100100111000101110100011001100000110001101011001101100011110001110111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out715[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out715, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110001101010111100111011011001010011101010101111111001111100101011010011101000001101100101101011101111110100010101101010110; 
out716 = 128'b00111000101110001100100001001000011001101010110000010011111101011110110001111000111010010110110110100110011010100001011000110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out716[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out716, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011000100101100010111100111111011100110111000110011000101100000010110100011101100111011011100110110100100100100110000111101; 
out717 = 128'b11101010100111000011011100010111001001111001100101011110101100101001001111100101110000011011010011101011101011111111101110111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out717[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out717, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101101001011000001010100101100100010111011101001110000111111110001110110001010010110111010000011110000011100100100011000001; 
out718 = 128'b01101000100110111000100000100011111001000011011111001101010111011101011000101001000101110001100000100011111111100111001011010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out718[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out718, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110110100010011010101100110100100000001110110001111010000011000101001101110100011100100101110111101110000111100111111010011; 
out719 = 128'b11100111100111010101101011101100000110100101010111011011100001101010100101110000000011101000011001110011110110001111000000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out719[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out719, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011101101001110100001101110110000010011100000010000101111001000001111100100100001101101010000001010101001111000110010001001; 
out720 = 128'b01010010100110011111110011111010010010001100010001000011111111111011001111001101101110111101101000001001011000101101001011001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out720[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out720, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111000111000101000010010011000000010100000011001100110101010011001010110111001001010010011010100010101111100100110001010110; 
out721 = 128'b10110101011000000010001101110010111100111001101111101011101001001000000101000100010111000101111110111100001110000001111011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out721[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out721, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100001010111000100000111010000101001110101001101110001011111001111111000001111110101001010101111011100110000110110101101100; 
out722 = 128'b10011100011010111001001011110101011010000111000100110111010001011011110001010110101110000101011101000110001111010010101000100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out722[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out722, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011110011101011011011000000000101011111011111101101000001101100111110101011001101101101100100001111111010010101001010110110; 
out723 = 128'b10010001001011011001100001111010000101101110100010111110111101100011110100001100000010011001110101111100010001110011100011100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out723[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out723, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111001000001101000010011101011010000010111111011000000000110001110111110110001000110010100111000001010110110110001100001010; 
out724 = 128'b00100011101111110001101111000001110001101011111001001100110000001101100010100100001011010010100111101011110100100110111011101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out724[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out724, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011010111001010101100010010100011100110010100101101100110100011010110001011100001110100100100101011100001011110000000000101110; 
out725 = 128'b00000010001100110110000101001001101100010001001101101000101010011011010011100011010111000101011000101100011110010100001110001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out725[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out725, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001101001000011100101100001101111100111011100101100101101111101101100000011000000111101110111100011001010001010010101000101; 
out726 = 128'b00100011000100111000111001101110111000101000011000100010001000000100110001100001111100001010001011001000010101010011000110011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out726[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out726, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110101101110111000101100010110110011101111011101001000001011001001101111001100100101111101110101101100011110111001010110011; 
out727 = 128'b01011000010001100011011101000010111100111000001100111110110001010111100101101010110000111011111110000100110101011001010001101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out727[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out727, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100101000001111101011000101111101101100011100011100110100001001101110111100010001010011111101101000110010101101101000101011; 
out728 = 128'b10100111110101000110010101111001011000010001110110100001111101011100010011011111101010000100000101111000011000010010101111001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out728[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out728, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011100110101111101100100010000001010000000010111110000111001001010000001001000011101110001101000100011110000001111111011010; 
out729 = 128'b01011001001000011011111100010011111000010010010010101101010100010100000100100101100111100010110010100111111111100110111110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out729[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out729, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001000110110101101110001101011111111111001000001110011001110000101110000110100110111001011001001111111000101010000110100001111; 
out730 = 128'b01011111101001011001000010100101001001010011101110110101111101101110011101111010001001111001001101010001001011101111001011001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out730[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out730, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011011001001011010100010000110110110000110011001100001101110111110000001010011001000110000001111001011111000011100010101011; 
out731 = 128'b01101111111001100100110010000110011110000010000100100100111001110100001110010111010010000000111101010011110000011111110101110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out731[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out731, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001000001000011110101101001001000010110100101010101101010100100110000110001111101010100110010010010000110000111110011101101; 
out732 = 128'b10110000010000101001111100000110001001000000100001111111100000111101101101011000101011001000110100001101010011110000011111001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out732[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out732, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001010001111011110000011001011101100100011101001010111010010110100011101110110011010001010110101110110110011111110101011000000; 
out733 = 128'b00010110001110010011000000110010111001000101101111010011100011001110101111110100101111100101111010001101111111010011110110001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out733[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out733, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000001001010111101110101000101100010000000000011001010010100110011000111010001111110100100100011001100011011110110101000111; 
out734 = 128'b11101011010110100110101010101110100100111001011000001011010101110000110000000001001100011001000000100111101110100111110110010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out734[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out734, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000001101111111001000111011110010100110011010111110111110111110010111101010010110100101000111100101000110011010100010111010; 
out735 = 128'b11010001001011011111010111010100011110110101101001101101001001111101111011010010101011101011000001010100110000111111001011000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out735[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out735, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111001011001001010011101100101010110010010011000101110110001101011000110100001110101010011010100000011001101110110111110111; 
out736 = 128'b10101101011011111101101000011101010111101100000001010000111110010000111101001010100100100111011000101110011111110001010100000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out736[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out736, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110101001000111001101010110111110000111010011110001001011010111000111100010000101110111001111100010000101111000001011010011; 
out737 = 128'b01000001011111101111101100101110100110101110101001011100101101111010111110000101111101110000100001101101110101010110101011011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out737[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out737, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100000001010010011110101111001101010011110100001110011001100011110101011100101101110101110100101001100101100010010000100101; 
out738 = 128'b01011101110001000010011100001010100110111101001010001110010101000001101000100101100010101010110100100001110001001111001101011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out738[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out738, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101110011101001010101010101001001000000110100000011100000000110100010000110000001110000000110000000101110110010000011000010; 
out739 = 128'b01001100110010011011100001000010110010011011010001110101010000010001110001011011100100001001111011010011001111001000001011011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out739[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out739, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111000011111111001011111011011111110111001010011000011100100110110111110111101001110010100101011111110111110101111011111001; 
out740 = 128'b00100011011001100000100111011010001011010110100001001101000010111011000101001101111000101101010110010000100100101010011001100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out740[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out740, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000110101100111001010011010111000111110101010110011111110101001100111101010111101110011110111100110011001011010111100101110; 
out741 = 128'b10001111001000011000011100001010101001111000010101010001110011001000001000111100000100101110100001101101100110110111000010111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out741[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out741, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111110101101001110101011001011101101001001110100100000101100010101001110100010101101101111110001011111101011100100011110011; 
out742 = 128'b11011001001110100101011001100001000110001010001011001000100101101101101110001110100100010000000000011110100010011000101010101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out742[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out742, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010101000001110110100010011011110100110110001010000111110010100010100100010001101110001111100011110100000010111000110011010; 
out743 = 128'b11100010011011110111011101111000101010110000000000011000111001101000100101011111001000101101100000011111000110101111111101010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out743[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out743, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100000011110011000110111111100001110001110001111101001110000100000000110010111101110000001000110100100111010111000010000001; 
out744 = 128'b10100110010010111110101011111000001100100100110110001001010111110100010000110000110101010100101011000010011100011001101100111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out744[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out744, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011010101100101001110000000111110011110111011001110010010010011100110011001111010011100111101000010011001101110010101111000111; 
out745 = 128'b01010001001000000100001011111100011111011110110100101110110011101110101011110001101110100000011100111110011001000011100100011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out745[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out745, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111011111111100111100001101011100110110011001100110110001100011110101001111000111111111110011000011111001000011101011100101; 
out746 = 128'b01100011011001100000111101111000000111101110101100010110111000101001111110010000001110000000101000100101110111010011110110111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out746[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out746, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110101010011000011001110011000001111011011111010110101110111111001001111111000110110011001000100101000100111111001110000011; 
out747 = 128'b00001001100111001010100111011110000110010000100110010011111010101011001111001011000001011000001010100101011101111010011010111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out747[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out747, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101111001011100110100100010011111011000010100100001100101010100010101001010110111110100001100111101110111010111111110000110; 
out748 = 128'b11110001010011010101010111101110100111000110100010010011101000110010100010001100101001000011000011100010110001101101001101100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out748[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out748, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100010001101000010101110111111100010000000110101101100000011101111101010100111001010110001100111010111110011100011011001011; 
out749 = 128'b01110000100100100110001101111101011010011001000000111010100100010010111110011111011010000011011111101100110011011100001111011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out749[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out749, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001111100111101100001001111110010011011110111101100111111001000100101100100000101011000111101010011010100000010010110000111; 
out750 = 128'b10110111101000011000110111011011010001010011011110011111000100010000110011100010001111100010000011010100011001010111110110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out750[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out750, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100111010110011001100110110100001101110001011111010000011101010101111101100011011011110100110100010000100100011000110010011; 
out751 = 128'b00000110111111111101001101001010000111111001000010011111111110111100001000000011100000100010110100011010010001101001111011001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out751[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out751, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100100000110100110111011110000111110001000110100000110111000101011000010011101101011101010111110011001000101010110111110101; 
out752 = 128'b01010011000011001101001101101110111010110111001101001111110110100010010001010111101011011001000110101000111010101101110000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out752[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out752, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011001110101011111001000101110001000001001011111101100110110001100110000000101010100011111001010001000111111011111011100010001; 
out753 = 128'b10100010111111100011000001101000111110011110111100111110101110000011111000111110101010100000101111101011111011100100101110001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out753[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out753, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011101110011111100010001110010101111011110111111011111010101100110110010111110000111111101010111011011110000111101010010100; 
out754 = 128'b00100001111000101111001101111011001110111011010100111011010001001111111001000001000000111111000010110101111001111111000101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out754[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out754, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100010000110111111010110001111010111000110111000100000100010001110011101001011101010100111110010011100000011010001111111011100; 
out755 = 128'b00110010100000110101011010001001111010100111111011011011000001010000011010011100101011100100001110100011011001100001010010011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out755[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out755, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110100101000101111111011100011000001101110010011111011010000100010010011011000011100000000100001010111111000001000001100101; 
out756 = 128'b10010111111100100001101100011100111000011000100110101001001100010110001001001111000110111111000000000001010001001111011011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out756[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out756, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101101111111100000011011101011100101110100011000110001010001100111100010000000101000110100111011101010110000011011100000111; 
out757 = 128'b10011100111011110011001000001010000101110011101010011101000110010111110110011100111000111010001001101010111100000101000011001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out757[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out757, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100101100101011001100100000110010111111100010010010000111010010000001110010001110100010010010100110110010010110100011000101000; 
out758 = 128'b00110100111110010101101000011101010011110000110111000010011110100000100001000101100000011100010100000111100010010110101011010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out758[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out758, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111101010101001110110101100000101001001110011001101001110100001011101011100011011101010011010101000100110010111011101000001100; 
out759 = 128'b00111110000101111110110000110000100001110110011000110001111000110010011111110111100100011111000110011110111111011001001010101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out759[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out759, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111000000100110110100101010111100010100011001111000011110010011100001000001101110111100011000111000011101011001111000101001; 
out760 = 128'b11101110010101100110010011111101001110111111001100100001111000000111011101110010000010101100000000010001001101111000110110011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out760[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out760, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101111000110011111100010110100010001111110100110000101001001101100111010010000101101100011110010111011110100111010010001100; 
out761 = 128'b10111011011011111010001010110001001010100111111001001011001000101111001011011000001101100100111011010101100010111000011111111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out761[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out761, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000010001011101011001010011100010000011101110110011001001001001011000000110110111000010010101011110011011110110110011110000; 
out762 = 128'b11001001001011000010101000001011001001010100101101001100100001110110011010100000001111000001011110100011010001101100010100111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out762[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out762, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000011001010101101000101100001010111011000010000001010110000001001111010011011101011100000101000110010110111110101111010110; 
out763 = 128'b10000110010111100100111100001011010110010000000111111011100000110100001111010111110110110000001011001001010100110110010101001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out763[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out763, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100111001011100001011000110000011011000100000000011101010011010001011111101110001111111000101000010101100000110011011001011; 
out764 = 128'b10011001001011000110000110111100100011111011100100011111110101010101011001010010011010100010001001001100110100011001101001011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out764[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out764, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110101111000101011111111000111000111110000010000101011001011100000100110100010101010100111001010001100000110101000110011010; 
out765 = 128'b10001000101101001111110101100010010111001011110010111010110111011111010111101010101011101001010101000001010010011111001100010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out765[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out765, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011111010011000011110100000011011001000100000000011101110101000000110111111110100010111000000101100111010110010100000110011; 
out766 = 128'b10011011011101110110100110110110000110000001011000111101010010101010001111101000001010110010001101101001110001101101011110110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out766[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out766, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111111001111110110110010101101000010111000000000001101100110010111101011111100011010000010010101101011000010101011100101101; 
out767 = 128'b10001001010100101100110010011011111011111100111010101001101110110001101000000000101111100110000000101000110101010010111010110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out767[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out767, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001100010100100010100100001001001110100110111011000010110010011001101010010000000111100000110101101000100001010001011101001; 
out768 = 128'b01100010010010101011111111101011101100101010100101100110001010001101000010100100101100011110100010001011111001001001100010110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out768[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out768, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101100100010011110000101011001111001110000011000000101000001111011011000001001010010000001010111010110001111110000101100110; 
out769 = 128'b01101101010000100100101100000100011110111010001001010001100000110010010111000101000000111010000011101110100001100011010000010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out769[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out769, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001100101010110010011001101100010001010000000011010101010010111111010010100000110011000111111010000111010110100010110010000; 
out770 = 128'b00010010100111111101100001001011011101001011101100001110101101011101110101000000101111100111010010100011111011011010111100011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out770[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out770, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001011000110110100011011111010001010111100001100110011010100011111011100100000000101001100011111100011101111001000100001111; 
out771 = 128'b01101100001010110100101100000111000111100011101011101011101000010101010111011101111111100111110100000000111101110100100110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out771[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out771, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101001110100101100001100011110001001010101001001001010110110000001111011011011110000010101100011100101100000110110110010011; 
out772 = 128'b00000111010110100110010011011011111110001100101100001100000001101010001011011110100000000000101001101000011111111111111101110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out772[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out772, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001010011111010111101000001101001000001101110101111001101011010101000000101111110101100110110010001111110010001101101010010110; 
out773 = 128'b11101001001011110101001010111111001011011111100111001110000100011011000110000000000100001110010010110000111001011001101101110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out773[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out773, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110101001010010001000001010110000001010011110001110000001000000000100011110110000001100101000010110001101011000011000000000; 
out774 = 128'b10101101101110000110100011010011110111010101101001110111110011001010101111000011001101110100001111111110110101011100100110100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out774[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out774, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101000101000101011000011001111111000010010111110111101011010110101100001101010010100101101001110111010011101110110010010010; 
out775 = 128'b11110110011100010111110110010110010010001100010110001001110110001010000001001111110000001001111010011001100110101111010011010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out775[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out775, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010110000100101001011100101010111101100101001100100000101000011011100000100110001101100111000110111000110110000001010111000; 
out776 = 128'b11111000010011000001011101100110110000101001110010111100011110011011001110011000011111000011000011000110101111100010111001000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out776[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out776, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001000010000011110100100010111000100100010001010000011001101001101011011110010011100111111001101000010101001110100011111100000; 
out777 = 128'b01010100100101101101110101100001011101110110010110101010100111000101011001101111010110011100011010101001101101010001110010100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out777[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out777, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000010010100010001000100111110101000000001110110010110000110000010000111110001010111110101110100011111101100000111011000111; 
out778 = 128'b11101000010100011001001001000011000100000001010000010011010111110011011101101011010101101000110110111101010100001001100000110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out778[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out778, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011001111111100001110001101000111011010111110011000010100000011101111100010000010100110000110010001001001111001100100011011; 
out779 = 128'b01000001101101001010000010100111110001000110010001010100100101010001000111100110110010101100010101100000010100111010111000111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out779[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out779, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110001100000000001000101111111111101010001101111000101010101001100101000111000110110101100100010101011101101001010101011001; 
out780 = 128'b00111000110010000110110101010110101011011110101010111111010110011111001010010001000010011010100101111111111100000101101001010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out780[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out780, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100001010010000011011000111101100011111001010010000000111110100110110100101001111010010001000000001010010110010010010011010110; 
out781 = 128'b01101000001000101000010001111001100111100000111010101010101111100111011011100110101110001010011001110000000001001011011100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out781[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out781, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110000101001001000011111111000001001110001111001100010001100100111001001010001110101110100100101000111000001110101100011011; 
out782 = 128'b10001010111010101011001110010110000011000110100110101110010110100111011000000111010000010011010001110010110110001110001000100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out782[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out782, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011001001001010111110101100011010000111101011011010100001111011101011110001000000011111101010001111010010010111110111110001; 
out783 = 128'b01010010111100011001000001011001101011011011000101110100110100111000111100000000010101001101011000100011000010010001111010011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out783[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out783, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010001010100110110100110000011001111001101010011000010100011110001100110111101010010100101100001100101101111110010110010110; 
out784 = 128'b11110100100001110100010001011000011101101111010010101111011111101000001000101101001011010010111100010101100000001110010110000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out784[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out784, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111111100001000011111000100000010110100010110010110110011110100100110001100011100101100001010011110001011110000001110000111; 
out785 = 128'b10101011000100100011111101000110000000001000110111001000101101010111101001101000010010101000101010111111111101010010100111100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out785[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out785, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001110000000010010110110101001010101010001001100110000011111011010111101011101011000101100101110011000100100000111010100000; 
out786 = 128'b00110011000001010001111100010111000011000110000110000111101011001110001101011000100001000111110011000001110111010000111100100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out786[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out786, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011011010001010100110001110101110111100001000100001111010010110111001100100100101011000001110111010011000100110110000100011; 
out787 = 128'b11110010011000100001100010101011000111111110100110011101111100010001001001110011110101011111111111010101100011100010000110011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out787[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out787, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110001111010111111001010011100000111110010001011111100111100000001001010101010100001100110010001110001101111100001100011001; 
out788 = 128'b11101000101000000011000000010110000100101101001110001000000001011000101110111110110100000110100001111011111100110110010011111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out788[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out788, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100011100001101110001000101000010101100010111000101011101111101010011001110010111100111101011010011000100001001110100000101; 
out789 = 128'b10001010000000000011010011011101001100000110100000100001011001010000011101111100000110100101111001100010011111100110000010011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out789[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out789, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111011001000100000111111101110010010111010001110111010011111100111100001010010001011011110000100110110111011111101111111010; 
out790 = 128'b01000001110011010111100101001011111010000111011100011000101001011110000110011101110010100110101000101010011111111011110111011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out790[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out790, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001110001111001010011110111001110110110111110000100001000010010001011110111011100101010100101001111011011100100010111111100101; 
out791 = 128'b10111110011000110010000100011000110110111000101000111110010111101111100100010000100100011110010000110101001000011011011011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out791[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out791, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000100010010000100001111100010010100011100000001010100011000000101111110001111010110111110010000101110100010000110111011010; 
out792 = 128'b10011000001010111101101000101011110110011110001011000101000010100110111110000111111000011001100110101110011001110001111001110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out792[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out792, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110110101101011100000110010000011000111110000000110110111111100100010100101100000011100001000110111001111101001011100100110; 
out793 = 128'b00001000111100101111101111101001101111111011010011011001010010000001001101110010011011000000010011100011100011011111000101011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out793[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out793, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111000000010011011001111001100001101010101001011100010001100100111101000000000111111001110011011000011010011101111111000111; 
out794 = 128'b00101110011011111101100001111001010010100100110101111110110100001111011000010011010100110110110111010111101101110010111001111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out794[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out794, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111101110101100100011010110100100000011000100111110011100001001111001111100101000111001010111101011101101001000011010101101; 
out795 = 128'b01100111011100011000101010001001111010110110011110010101010101001000100011010010001010100000101010110000000111111000001011001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out795[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out795, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111111000010101110111010101100111111101001001100111010100100111011110001010011010001011011110111010101100010111001001110001; 
out796 = 128'b00111100000001111100111100101011000001000111100111001010110110101001001010000100010010011011101011111011000000011001101111011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out796[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out796, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111000110100011010101010111000010001100111000000100000011010001101011100011001111000011100100001111010000000001011111101011101; 
out797 = 128'b11101010011110001010110000000011101111001100101001101110101001110010001110011011011110000111000100111011100010010011100011111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out797[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out797, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100101011011110001101000010111101101010100101100010110111101110101111011101111100000100111110000101100001111110110110011001; 
out798 = 128'b01111010001010011000100010101010100101000111101001100011100010100010000000001101101111011000001010100000000011101011100101100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out798[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out798, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110001100001001101111110100110001011010001101011101111001100010100100010000111011010010011101101100101111110011101011001101; 
out799 = 128'b00001010011100011010000011110010111111001100000100111001001101001001011101010000111101000001011111100001010100101010100001000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out799[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out799, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111110000011010111101111000000001010101110100100100111011010011111010001010100011101001101110111111010000001110010001100010000; 
out800 = 128'b10110110000011010111010110011001101110100000010011000100000000111001111100110110100111011010110000011010010111100110010100111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out800[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out800, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101101101111111001000010011001111111111001110111000110101100101001111111000001111111010001011011101010101110110110000110110; 
out801 = 128'b01011000110011010100011100110100000101000111100011111111001100111011110110111110010011111010100111010010000111011101001101110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out801[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out801, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001100000101111110010110101110111000011001000110100010001100111101000000100101100111001110100000011111011001101100100101001100; 
out802 = 128'b10111000101101100110111000101111100110110101110000110010010001110010010100011001101100101000011000011011001000001111111110100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out802[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out802, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000010100001100101010110110001000100011111101110011111011101100011011111011100101010100000010101110101110111111111100010101011; 
out803 = 128'b10110110000000101110101001100001011101011100001110010010011100110100000001000111110100001000100000011110011100000111010000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out803[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out803, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110110001011010010000101101110011011101111001100110010111111110000111001110010001000001010000111110100001100111110010010110; 
out804 = 128'b00000110001001101101100010011111100010010001100001000001001001001101100001100110010001010111010010001101110100010110111010001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out804[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out804, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111101101000000001001100011110011000100100001010000011100000010100000011010010111000111100110101111000001011000100100101110; 
out805 = 128'b10001100001000101110010100111011101110010000010011111011110011000001100110001100001110101110110110101110001011001010100100001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out805[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out805, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110111101001000010001011011000011110100000110101100000111101100101110110000101111001101001111001010010110101111001110010011; 
out806 = 128'b10101000000001000001010001110000100111010101101101100110111100011101010011011010010111011101000010001001111000010111101100100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out806[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out806, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011000100010111111011100101010001111110001110000000110010010010110000100011011000111011110011110110110010110000101100000100; 
out807 = 128'b10111001111100000111011100000100010011100110101001011110011101110111000110100111100010001010011101111111011000101110101010011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out807[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out807, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101011000011010010100011111011001010011111100101100111110000000111010001010010011101111000111101101110011111011011111110100; 
out808 = 128'b00010111011110010101110000100010101010111110100010110111101101010001110101011010000000010110111010100000110000110001110111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out808[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out808, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111101100000101011010000010101010001101001111000110010100111010100000001110101010001000001000010110111110000111110010110000; 
out809 = 128'b11101010011010111011000111100011010111000000001010000101110101000011100000011011001001110110001001100000000101101001110100000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out809[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out809, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110100001000101100010000000101101011010001001101010100100001010010001000110101110010011100010011111011010110100111100111100; 
out810 = 128'b01000010000110000010111100101011001100010111111010111001011000101011111110101010001100001110011011111010001100001011011111010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out810[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out810, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111001010110001110001110000010000110010101001101101010100100110010000011011101011111001100111100100101000000011010010110000010; 
out811 = 128'b01110111000110001000010110111100110011101110111110110011000111010000100101100010010000000000101001101111000011000010111000010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out811[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out811, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001010110101011010101101111111000101101111101001101011010011111101011010101011110111101101110111110111111111001110000011000; 
out812 = 128'b10010111110011110110101100001010111011110100000111010010011110011111000111001101100111101001001001010100111010110000000001001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out812[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out812, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111111001011100001011110010001000001011000111011011110101110001111000000111000110100111111100011010110100101000100101010000; 
out813 = 128'b00011101111111011100000100111111011011100001100101101101110000111110000010110111101001000011001100010100011000101110100111100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out813[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out813, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010010011101111000001000001001000111011000111001000000101001100011000111110101101100001001101001111110010010000101101000111; 
out814 = 128'b10100001100101011110010111101110100000000101000001110110001001000111111101001100011100001011001111100011111101001110010011001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out814[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out814, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100101011011100100111100011101010010111000000010010110001110011110000111010010111110100110000000101001100110100101011100010010; 
out815 = 128'b00100101011111111010011000010100110100011011000001001101001000001000110101011111011010010001010110100110000111101110000001111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out815[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out815, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111110110011011011110101101010100100111100001100010111001101110101100100000100100011110111001110110110010010101111110110011; 
out816 = 128'b11000011000110110110010010001100100000010100000111101001011001000110011101110110111110110000001100100111111101110000010100101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out816[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out816, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001100011010011001110000111010111110100111101011011100100000110111101001101010001101010110111101101001001000110100011100010; 
out817 = 128'b00111100100100101100101011110111001001100100011111011101011101001011110011001001011010111010001111100111010111111110101110000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out817[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out817, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011111011110001111110100010010011010011101100000010000100011110100000000000000110000010111100110101010101000100000110100110; 
out818 = 128'b01000110110010011110001110010111011000100111001100010000101110011110000110011000001011001100000010001101010101001011010001011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out818[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out818, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001111010010010110110000110110000100110000001110111111010101110111110111011100110111100010101011110111010001101001101110011110; 
out819 = 128'b00100101010110000000101011001011111110010000100100001001000111010000101000101011011110100100101110010100101010111100000000001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out819[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out819, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100100011010101000011110100010100010001011001100010100000000010011100011010000100100010011100011000011110000110001011100100; 
out820 = 128'b01011110101100010111001111101110110101100001011101010001100110001100110111110011011011110010101111101111101001101101110011001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out820[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out820, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011100111010100011010101000010001100101011110000110010011001100111001111000001000010010101111010011000011011100011100010010; 
out821 = 128'b11001011100111011111101101100100101100011111001001111111111001000101000010110000111111101101100001100011001110011001010011101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out821[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out821, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010000110110110110101010111100000100100111110011110010101100010101000000011110011011110011010000001001101111000011010001001; 
out822 = 128'b00100010010110100010001001100111111000001100000010001001100111000101010100000001100000110000010010010001000001010010110010011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out822[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out822, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010010001110011110001101001110111110010011011111011110100110001011111100010011001111000000110110101100010010101101001011000; 
out823 = 128'b10011110000110100010111101011011100000011110101111101101100000100001110010101010001100100011111000000010100101010100100111011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out823[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out823, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000001111100110100110101010011010101111101010101011001010001101000100101001101011000010111010010010111111001001011101101101; 
out824 = 128'b11010101001110010000100100011101011000011010000000010111000100001011110000101101011001000010111111110100011111011110110010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out824[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out824, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100111010001110000101111000110110100111001010110001001111011110001101110111100110111101110001111101010110100000001101110011; 
out825 = 128'b11111000111101110001001100011010110000111011100100110110111110100010111000110000100101010000111101011110110100110010101100110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out825[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out825, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101011111001101000111001000011110101100001101000111101110011010100010011001011111010111110001010001110010000011011110000101000; 
out826 = 128'b10100111101110111001001000111111010101010111101111101011011101111101011110010100011110001110110101110010100110011001101011100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out826[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out826, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001110000010101000000000111100001000101101001110001010110111111001101010010010000001010100111111011010010001000011001100101010; 
out827 = 128'b10001100011011011110100101001011001010110011001110001010100101010010111011111101000000010000000111111001000100001011010001000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out827[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out827, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110101010111111001011011000011111001000001110100001110000010010011001011110000110110101111101001111101001010100100011110001; 
out828 = 128'b11010101011000111000101001110101011111100000000011111111101101001011000001110100110011101011101001010100111100011100110000010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out828[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out828, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011001111000111111101010101101100111010111101110011100110111111111000001101101001111000011111110000001011011101001001111000; 
out829 = 128'b01101110000001000100101000001111111010001100001101000010010010011000010000010100001000111000001000000010000010010010110110010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out829[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out829, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010000001010011000011101000100101011110000101101100101111000010011010011001001001110010111010111010110000111010101000111101; 
out830 = 128'b00001010111001110100000011001110110011011101001011010100100010010101111100111001001000101011011111011011100100100000101011010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out830[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out830, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010000101101100101001011111001111110100111110001000000010000101000101010111101100000101000000100100000111100110011110010010; 
out831 = 128'b10111110010111000010001101001100111011101000011101100000100001101111011100101000001011000000010011110010000101000111110111001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out831[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out831, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010111100101110110011110010110001100110000111100011010001111011100101001000111110010110001101111111010100011000101101000000; 
out832 = 128'b11110000000011001011001010001100011000100111001100111110111010010110100001010011111111111001001011111000000001001000011101010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out832[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out832, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011111111101110010001001010011100111110011101011101000100011000111101011001010000010100010011111010011110001011000010101001; 
out833 = 128'b01110001111000001101100110010100001001111110110111011011010011100111110111000001101001110100010000011111001110011001111100000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out833[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out833, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000110110000101100000110001101111000011001000000000100010010101101100111110011000010100001100001010011001010011010011111010; 
out834 = 128'b11101111100101001011100000000100100111000101100001100100010101101011010101100111100011010111111000111111000110010101110100000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out834[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out834, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111011100100101001010011010011000000111011011000111010110010110010001011010001110001111010100100101000101011000101100011010; 
out835 = 128'b00010011101001011111011010010001010111010110111011110010101010101111001100101100011000111001100000100000000001111101011011001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out835[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out835, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000101110101001000101111000010000111010000111101010001011100101100110011101010000101000101111011110111000101110000000101100; 
out836 = 128'b11000011001011011000010111111101000001110110011010010010101010011001111000010100111110111100110110110110100001100111110100010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out836[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out836, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111011111011111111110000110101011001001111011000110111000001101101111110110101010001111001000100010110000100000001011011011; 
out837 = 128'b11010111101010101101010101110001101110110100000100100011111001100100000010011101110110110000111110111100101100100010000110111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out837[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out837, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100000011111011101010001100000110001010010101111010010111101110101101000001110100011011110101000100100111111101000111110010011; 
out838 = 128'b00011100010101010011110000011100010000100000101110111001100000011110010011111011000100001100100111111110011100000101100000010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out838[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out838, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010101001010011000001100110001000101011101111001101111010011010110000001110000110000101111001000110000011111001011010100111; 
out839 = 128'b01110101111011011001010011001101101000001111010110110100010010101000101101111101101011010101101001101001101010001001100011110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out839[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out839, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111001001111101100100000100011000110010010111100111110001101111111111011011000001001101011000111110010000100111101111000000; 
out840 = 128'b11010111110001111101001100101000111000011001001101001111001111011001111000100011100000100011001101111101011011101011101100101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out840[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out840, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000010001101000110110111101001111001111110100110101110010001011010010000001101011000100010011110111101101010000100100010000; 
out841 = 128'b10000001110110100010111000001011111101110100011001101000101001111100001001010101101001001100111011111101001000110010011010011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out841[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out841, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110001010100110100001010011100100001111011111101010001010001101100010000000111111010110001101010100100100110111100010101100; 
out842 = 128'b11101011100011010011000111011110100110011001010100011111110101000001001010111011010000110000111001010001010100100111111111000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out842[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out842, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011011001110001000011010100100100010000111100101100101100100000110000100011111110000000101011011000111111110001011110011111; 
out843 = 128'b00111001100000110011100101110110111000111000000011000001000011110000111111001100111011101010110001000001101100111011000001000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out843[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out843, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100000101000010001100010000100110001111000010100101011010000100010010111010000101010100000101011111000101011101101001111110111; 
out844 = 128'b00111000010010111011001110111010111101001110000011010101001110000010110101001111101100000110010110101100111000100011011001011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out844[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out844, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000010011001111001001110111110010110000101101011101010001011110100010000011110110100111001000001001100101100110101110111001; 
out845 = 128'b10101100111000101100011110100100100100001101101100011010000100100111001101011000011010011110100000001010101011001100001111100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out845[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out845, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101110000001111000010100000011110011011111000101100010110111101010001000000001100100011000110100111101000110110010000100001; 
out846 = 128'b10011101010011111101111001010000000011100011000010101001100100101101011100011001111110111110110011010011000101000101110111010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out846[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out846, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010000110110001111111000011101111001101000011100111001000011000111000010001101111111010001000001010101010111101111001110001; 
out847 = 128'b01000101101000101100000010000001011111000001010101010000101101110010000001000101011110000110111011010010110000101101100100110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out847[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out847, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111000111001111010100100000111100110001010010100100010001110110100010001111110001001000011000111000111000101110110101111001; 
out848 = 128'b00100010111010011011100011111101010111110100100010001110100011110111100010011011011011101110100100010101011011111110100011100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out848[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out848, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011100101011010001100000011110111000000011001111101111001111001100111001000100010101000100100010111010010100010001001000000; 
out849 = 128'b00101110110001101110000011011010001000110110101110111110001011000010010001111101000000010011001100101000000101101110010000100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out849[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out849, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011110011011000110010010010010111011111101111011110101010010001101100100101101010100001001100111111101101000110100011010000; 
out850 = 128'b10000011101000110000101100100110011001000010111111010001011111000111101101011010010111110110110101000100110101010111000110100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out850[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out850, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010010000011101000001110111010111101011000010001010111110000011101001000111010000001101000000101010000110011110101010011010; 
out851 = 128'b11011011000000010111110110101100111001000111010000110100000000011100101000110101111000000001010110000100000000011010001110111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out851[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out851, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110011100111101011011001110001001010000001101011101111111101110001111010100100101010111011000110110101101101011110000010010; 
out852 = 128'b01010000101000101100011000100001101110110110001100101000100001101010011001010101011100010000100000001111111010110101100110001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out852[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out852, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100001001100010001111111010001001110011000000001101011010111100011100011010101000001000011011101011111000100010001101011010; 
out853 = 128'b10001000101110110100111000010011111110101000001001110111111010001011101000111110110111110101101010110011001011111100101011110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out853[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out853, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010111110000001011101101000001011010001000100110100010011011010010110000001010010100001100010010111110011101010101111000011; 
out854 = 128'b01111110001110111000001111110011000001001000110101001110000010110110111000111000011100100010111001110011011101011100101100000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out854[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out854, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111000100010001100111011000001111000010001110011010100101111010111010010110010000011100000011000110111000000101010111011000; 
out855 = 128'b00101011010011110100110111111100010101110111011001101110110010011011100010111100001011010011100001011100110110011000110111000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out855[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out855, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111110011111110101010000111010100110011100100001101111100110111110010100010111011100110100011010000011001010011110100100101; 
out856 = 128'b01100101001001101100011011001110011110010111001100100100111010010100001111111011101111000000011000100010110111111001101010111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out856[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out856, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111100001101001011011001001011000111010000111110101111111111101101110100101111111000011001001001100111000010011010101001101; 
out857 = 128'b00011111111011000001111001010101011111010110111010001101000001101100111100101111010101111011110100010001000010100101010110011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out857[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out857, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001001001000100001011111100001110011011010110010011101011000000100010000101100001010111000001100101000111010111010101000010111; 
out858 = 128'b01000101010111100100011011111010111011010000000101011101001011001111110111010011011011101101111101100101010010000001011100100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out858[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out858, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101111011111110111111010100110010010100100001010101101001000000010100101011111110010110110000110010110010101111110001000011; 
out859 = 128'b10010100010011000111100110100000111000011000110011011011000010111100001100001011100000010111000100011011100111110011101000110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out859[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out859, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001100100000100100011111110100101001110010110001100000111001111010110010110000110100100000001010010101111101100100011001000010; 
out860 = 128'b00011100111101000101011001011110101000100011011000111011010000101000000110010011100111011000101011001101111001101011001101011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out860[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out860, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011000001100110010010111000010110001101011100001001100110000000100001010000100001010000110000111101100001011101010110001111; 
out861 = 128'b00100111011011010101100110100000001010100100101000010001010000100111100100110111010101110001111011001010010010111010001011010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out861[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out861, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101110010110111111010111110010100101111111101000001100101011000000111000011110111100110110110110010000010100110111001010000; 
out862 = 128'b10000000110010010000111011101000001110000110111110011011110011101011101001101101000000100110010100000111000101111111110100110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out862[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out862, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010111100101111100111111010110101000111110101110110110101110010100010001000110111110000001000010001001110110110010010110100; 
out863 = 128'b11001011000011100100010100100110110100001011010111110101001001001011111010101100010011001100111001011100101000111100001101011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out863[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out863, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101100000110011110100111001011000001010110011101011010110001110101101001100001110000100011000101100101110011000101110100010; 
out864 = 128'b01000110110011100000100101111010010101101011001101001101110110010111011110001001000011010001001011000110101010000110011100111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out864[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out864, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000001011011100001100001100111001101000110010111000000011010010011000010111101111100010111110011101000100011000100101111101; 
out865 = 128'b00001110010101000000110011010000000111101001101100000100001111001001101001111001010011101111101010001001110011010110101101001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out865[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out865, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110111000100010100111010100111110011010110110010000111000111110110111000010001110011111011111011001000110010000011100100000; 
out866 = 128'b11101101101110010000110000100000101100000000000111010010000111001100011011010011001100100110100010100011000000110010110100100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out866[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out866, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101000100010000010001110111000000000000001101111100101011100011111010101010001110110100101101110000111011000001101101110000; 
out867 = 128'b11010010101101101010010111000010000000111000111001111001010111010100010000010001111011010111110001101001010011010000111101101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out867[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out867, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101010011110111111110010010111101000101010110011000001010110100011101010011100110110110111001100001010111000100011010011000; 
out868 = 128'b11000101001110000000100100000001011101010010100101101010000110011110110110000001010100010100001001100000000110001111101000010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out868[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out868, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101110110111110000111111001100100111110100000101011000000010101100100001110101100011111000101010101110101011111001001000101; 
out869 = 128'b00000001011001000110010110100100000111000101010101111101101111010010100011001101110000100011011010100111000111000110100110100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out869[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out869, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010010011100010000111011100011001011010011101010101001001100011011011100011101110011011110101101111111001110000010001111000; 
out870 = 128'b10111010011100010101110011011111110101101010011101000101110100110111111000111100010010011001001111011010101101100001101101011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out870[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out870, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001011100001010001011011001101011010110000001100100000100000001010010101101101010100001000001110011111001000001001111010111; 
out871 = 128'b00000101101110000001110001011000001100111110100110000001101101110111100001001100000101000000010100110000100011001111011100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out871[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out871, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111010100101011011100011101011011001001011111011100101101001111111100000110100110100011000001010000010100011110010101011111; 
out872 = 128'b01111011011100110111000101000101010111100000011010001111001000101000000100100010101011001000000001101000100111001000001111110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out872[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out872, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011111001101000010101000010111001111001011011001000001111111101011011101000010101100000001111101100011000001111100010101101; 
out873 = 128'b01011011000100110010110010101010100011000010110001100110011001011100000100111110011100011110011000010100110100110011110100000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out873[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out873, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111000111101101001001101111011101100100000010110000011110001100000010110010010100010100001001100110010111010011101111100001; 
out874 = 128'b11001011101010010111001000101000111001101000111111011011000101110010111100110110000110001010111011100110001101010000010111101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out874[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out874, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101011111011000000111010001111111101110010100001001000010010101110000000101110101111010100100100011011011010111100001110010; 
out875 = 128'b11111000101001100110010111011000000110111001110000001000000011010010011111110011000110110110001011001110010011110101100000110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out875[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out875, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010010101000110011010001011011100011010000100010110011001111010010011010110001000000011111111101011011010010000101011111101; 
out876 = 128'b11001001111001101010001110001010100000011011110100101001011011011100010001010100000101010101001010111111011111111001001011100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out876[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out876, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000011010010110011110010100001011010000100111111000001100010111001000001110101011101011001010001011010000010110010110010111111; 
out877 = 128'b00011011100101110111110010010101111100001110100100001011000111010001000011011000011110010111010100110100111010110100110000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out877[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out877, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100001110011111110001010111111111010001001010001001010010011100001111010000101000001011101000101011000010010011000010010010; 
out878 = 128'b01101001111101110100110111110001101001100110110110001111001111000011010011011011111110011010000001000011100110101111001010111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out878[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out878, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001101110010100101010100010011011000101000011010110011010100010100001111011110111010001010001110001001101101110101111000101; 
out879 = 128'b00000000010001111001001111101011101001011101010001011001111101000110001101010010000100011001001001011111000101110001001110110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out879[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out879, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001011110100110011100111100111010000010000011000100010110100000111000101000100000111101001011101111000011000000001110000010111; 
out880 = 128'b11010101110001010001101110110011001001110010000111110100101011100111110110100111001000010111010001001101011010001111011010111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out880[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out880, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011101000011000010000011011001111110110101111011010110110000110101011011010111111101110000010101011010000111100010011110101; 
out881 = 128'b10011010111101010011100011111101001011010000101011011010011110011111100110001100000110111111010010100101101101111011111111110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out881[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out881, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111101110110110101011001101111001000101001111111000001000011010000010110011001110001000101000011000101000010110100011111000; 
out882 = 128'b10000001110001111110100110010111100101001100101111000110001011000000000101111001110010001101000000111100000000011000011001111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out882[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out882, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100000001011100011011110001010110110001010001010101101111011101101101011011100110000110110111100101000101001100110101001100; 
out883 = 128'b00100010011010000000010010010001011000111010100001010100011001010100010000100111000000001100110101110100110010001001011001001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out883[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out883, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011000111101001011010101001101000100011011000101001100000001101010110110101001001011000000110010111010100011010001000000100; 
out884 = 128'b11001010001001010011101111101110010101000010110101010101011111000000001011000000010001001110010000100110110101000000101011100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out884[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out884, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001010100110001101101001011010000110000011110101010000001000000101010011011111100001111001100111111001001000000011000110110100; 
out885 = 128'b11000111110001110100101111100001010110011111000101100010111011001101100101000001000101000011101110100001010111110111000010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out885[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out885, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001010001001101010010110101010110011001000001111010110010000001101111100101000000001001110010111011110100101011111101100100011; 
out886 = 128'b11111011100010110111110011100010110001011100101000000111000010110100001011010101011000110110011111010010101000000111011101010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out886[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out886, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011000011000100001011010010010001110110000101011111110110100010000011100101011000111001011000010111100001001100111101111001; 
out887 = 128'b01000110010001111100111111111011111111010110001111110111101001011100110110100000011000001001010001001110001001010101010010100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out887[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out887, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110000011011000010100101101010110111110101001101111110001101011111000010011110011111010001001000001000111000110101101001100010; 
out888 = 128'b00110110011010110100011111101011100101111011101100011111100111100011001010101110101010101010111110001000100010011000000011110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out888[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out888, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110011110111100010111001111111010111000010100011111111011100100011100110001011111000010101101101100110001111011111110000000; 
out889 = 128'b00101000111110101001111001011011011001100000101011110101001011000111111101101010110110110101110101111100000000100100100111011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out889[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out889, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010001101111000100000000000010101010110101010000111101011011011000001101011110011110100110101110000011111101101011011111011; 
out890 = 128'b01011010100001110001010001010010110010110001100101111000001000001011010110011000010101100101100110001010010110001101100100001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out890[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out890, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010000001110010110101110111001001011101111011100111010000110101010111011100101010000111010010000111011001100111000001100111; 
out891 = 128'b11011110010011001011110110000010100100100000111110001111000111000011001101011110111101100111110100000011001010000001101111110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out891[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out891, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110110011101101011000011000000000110011100010101010111011011010101110110111110111010001011011111100000011101111010100100100; 
out892 = 128'b10000000000100100110100111110101100110010001110001010110101100111111011001001101011010111110101101110111011011101001111110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out892[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out892, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010000000110110100011001110011111010100110101001111011100010101110111110101010110111101110111000001001100000110100001001111; 
out893 = 128'b11011001000111101111011000000110000110111010000100010001101111010010010100101001101000001011111000011001110111100001100011001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out893[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out893, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111110011101100111010100101010001000101010000111000111011101000010010000001001100110000100000000000010010100011100100010110; 
out894 = 128'b00100011011000011110110100100100000011101000100110111110010100001110001100000110001101110100010000100101111000001101101001001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out894[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out894, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110011100000100110010110011111000000101101000101010111101011011100101011101011000011100101010110010001111101111110100111100; 
out895 = 128'b01010111000100000000000110100010001110110111100011100110100110110111011001101011101100011100111001001101010000010000101000001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out895[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out895, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010000101000110011000011100000111111101111001010000010011110100000011100000000010110111111111100100111000001000100100000111; 
out896 = 128'b11110011101011100011011011100110011110001001011101001000010110011101111010111100101100010010001111101000100100111100101000011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out896[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out896, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110000000110010010111000010101010110000000101011000101111000101100111001001111000100110110000010110011001000110111000011011; 
out897 = 128'b00000110000011011110111011110101011011111101000001011111100011100100110001110010001101000111011001111101101100111101101101001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out897[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out897, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010011001011000111010011000111011110000100011000100001000000000001010110001111100010010100111000010101001001001000011100010110; 
out898 = 128'b10101101111010100110100001011010001001001001001100100110111111100000000000011110110111000001010101111010111011100010000000010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out898[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out898, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000100001111010000100100110011111100011001000011000101011100001111110100111111010111101111001101000101011110111100101100110; 
out899 = 128'b10100100011011010101001100110010110001100100110111110100000111010010001110000001111000110000001111011011100101111101110100010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out899[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out899, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101000111000100110110000011010001011100110011010100010000110011000110001011001001010111110001011111010110000101011011001101; 
out900 = 128'b10100101001111010001101000010011100000110000111011111111110010100100010110101100101011011110101000001100001011010110101101111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out900[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out900, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001010001101111100000100111100001011110111010000001000100111010000001111100110000110100000001100111101101001100000011001010; 
out901 = 128'b11000110001110000011101010101011101100101001010011010001101010011101101011011110100011011100100010011101101001111101110010100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out901[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out901, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011110110110110101101011101101010010101111101011011011101111000011000001100101000011000010110010101000101110010001111001111; 
out902 = 128'b11100000010011010110001100001101100111011001100101101001101010011100010111100110001011000101110010010001000000110101100101110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out902[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out902, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110111011111100000010101001010101010101110011110111100001111010111111001010011100011100110000101011000010101001011101111001; 
out903 = 128'b01111010010001100010010100111100111100001101011000110010111010111000001110110100111010010100110111111010010111110000010000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out903[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out903, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001011001001110011011000111100011010111000000100000001010000110010001010011101011100010001000001110110110101100111000011010; 
out904 = 128'b11100000100101010110011010100001111010001110000000010111111110110100010011001001001010000011101101101100011000010101000100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out904[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out904, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011101111100111011000110110001001000111000001000100110001100001101110100010111111011011101101011001100011110101010001000110; 
out905 = 128'b11011110000101010000000111101101110110101100001101100111100111010100101010000101110010111110010110001111010000010011100000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out905[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out905, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100010001101100111100000101011010101111111010000010001001110001101011011111010010100110101101101101000110101100001111111001; 
out906 = 128'b10110100000001001110110110010110101001011100111000111010110110001110011110011001100001000010000110101010001000011011100100110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out906[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out906, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111000101000001100100101010001001001111110101101110001010010110011100000110001000110010000001101010010011010101011111011100; 
out907 = 128'b01100101000110010000000111001101010111110001111010110011011011010011111011110000001001010000001010110100111111100111000111111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out907[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out907, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110100000001101000100011101000100101100011010011100011001111111100011000000100110100100101001100000110101000000000000011010; 
out908 = 128'b01111100111011111100111010000101011010111101100000110100110001001010100110010100110010100100101110100010001110101010101000110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out908[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out908, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110111001100000110011101001001001100111001010001101001011110101110011000011111011011110110100000100010001011011100000111110; 
out909 = 128'b11010000011111110010101101010001100100011000011101100011001011111001010111011111111001010111111011100100010101001010000100111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out909[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out909, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011100010111101000101101010100010001111010011000011000001101011100100011100011000000110111110010111101111001011001011001000; 
out910 = 128'b00100001010001111001000010100111000010101010100110111100111111010111111010100110001111101000011100111101110100111101010011000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out910[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out910, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000110100110000011000010001010001110100001010011111100110101001000010111110111010100111110101000001000110100001101101000010; 
out911 = 128'b00111001011110010110101010000101111111100011001110000010000111110010000011000010000101000100000010001010011111100101001000100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out911[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out911, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110000101101011001001000110010101111001110101100000100111001010000110010110000000101010111100011100000001111101000100000101001; 
out912 = 128'b01010110001110000100100010111011110011100010011110110001101010101101111011011100100100011100111101110010011010111011000111100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out912[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out912, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011011011101110111001000001000111101000111111101010001010001110111100101000000011011001111111100010101111110010010100010101; 
out913 = 128'b01111110010101000110000111100110011010011000001001101100010100011101011110000000000110010111010011000110001100111100100001001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out913[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out913, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100011010000001110001010011010000011101000100111110100011111111100010110011011011001000001001010101100101010100001101011111; 
out914 = 128'b10011101100001101101000011111001111010011011011001110011101010011000000010000100001000010010010010001101011101110001111011101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out914[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out914, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111001001010100000100001000110001101001011110111001010111100101000100100001110011101011011000101001100100010011000001101010; 
out915 = 128'b00010001001100001010001111010110100111001001001110010010100000101111000010001011100011010111111001011010001000101100101010100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out915[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out915, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011111111001011011011011011101010110101001010100011100111111100010001111011110101110111011110110101111001010100000011001011; 
out916 = 128'b11111000100010000110100001010110010010000100011011010110001110000010110011110110101001010011000111001100110011001001100011001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out916[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out916, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101101001111001011110000101111000010100110001011101110111010010001001101000111111111010101001110000101100111100110011100011; 
out917 = 128'b11100100110111010010101000011011111110111110000000000101100110110000100011110110111110101100110111011011001111111011001101011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out917[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out917, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000011011000010111100111001001101101100001011000010010110001011010110000011010100100101110111001111111000100010100101100111; 
out918 = 128'b00111010111010101111111000010010001101010110001011111000101010111010001000111001101010011011000010010011011010111101011011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out918[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out918, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111111000011111011111010100011000010011010100001111111011000101001010100101110011000110110100110001101001110101000111011100; 
out919 = 128'b00011100001111111101111101011111011001000111000011000010111011111111100111100111101101000111010011110101011100110101001100110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out919[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out919, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001101010101011010001010110111101100001111100001011001010101101100111101100111111110101111100001100101001110001101000010011; 
out920 = 128'b01010011000001011110100111100100100001110011011101011110001111100110101011010000100010001010100010001100100101001001011111111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out920[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out920, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111111010110010001001111100111011010000110110110011011000011100010000000101000011110101001001101101000101011010000000000000; 
out921 = 128'b00110010111011011101100110100101011000100000101100100000110110000001100111010100010111010101101100000011000100111010101110010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out921[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out921, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001011101001101101000100011101011101000010001100001010110000111001100101110011110000000101010110001001100001111100110011010110; 
out922 = 128'b01000101111111000111110010001110100111100100110101100011010100110001100111000101111110111011001110101011011100100110101000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out922[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out922, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001011001001011010111011001000010101001011110111110010010011111110000000010111100001100100011101100100101000010111011100000; 
out923 = 128'b10001100010000000101000011000000100000110101100011010011111001111111011000111011111010000011101010011010100111110001000000011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out923[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out923, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111101000001011100011101110100001001000111001111110101111001011100111010010111001001101001100101010001110010100000101110110; 
out924 = 128'b00111000001000011011110111111111111001110100001010001000110100001000010101101100001110000001011011000010100100111101110001101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out924[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out924, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110110111001001011001110000001011011010111110100111010001101100110101010111100011011000010101000110101011011101010101110111; 
out925 = 128'b00100110111010010000110001010111110000000000001111000000111010100100011101010110110001000110010011111000001010000001011011001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out925[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out925, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011111100011100100100001100111111011110001001001110010010000100000110110001100100111110010111001100100001011100010001101000111; 
out926 = 128'b11010111110011011101101110100010111100011111100001011111111010001001111010010001010100110011011001000001010100101010101110111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out926[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out926, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010101110110100011000111110100001110111011000001101010001101100000110011010100000011011000011011001100010010011010000000011; 
out927 = 128'b01111000111101101010100001011001001001010110110010100010011111101011000110010000100010100000101010010110011100111000101010111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out927[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out927, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011110010111011010000000011010010110010101010001000000111011100101101000111111100000101010000101010100101110010001000001001; 
out928 = 128'b10111000011001001111100100110000100011000001100101110010011110111001110101001111110101000000111000010010011000001110110001101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out928[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out928, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110000000000010011001010111111000100101010110111010100001110000010100000011011100000010001110110011010001111011010001011111; 
out929 = 128'b11010000100010100101101001000101010101001001110111001010111111110011000100100111110101101010100000011011011111000010001001010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out929[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out929, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110011101010011011100001011111100110000011001110010101010000010011011010111110011100111001011100010111010010001100111010011101; 
out930 = 128'b11101100111101001010101110100110001110001101001111100001010111010100000001001101001101110110001101110000110110101101001000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out930[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out930, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010011110010101111110100111110000001011101101111111111010011101000000011111010100000101010111011011100100010001100011111011; 
out931 = 128'b10101010000100100011011000101101111111010101001101101100110001010011011011001000000011100010001001001011010001100011011101110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out931[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out931, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010110111110000110010011001101111001011111100110010000001011000100001010010101011001100110110111111000100110101101110001010; 
out932 = 128'b10100000101001111001101011000000100100110100001100111111110000001001000101000110011000110000010010011000000010011000101101110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out932[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out932, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001000111110111011110101111001111111010111101101000010000101110101011100100011000100000000100011011001111111011011000010000; 
out933 = 128'b00101001000111011110000100111001011111100100110101111100000011100111000001001001110011010001111101000111000101100100101000110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out933[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out933, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010110101001011111110111110010000010010101101011100010110100110111101001001110111100001100011111001110111101011110101100100; 
out934 = 128'b10011001000001111110110011100011011010000100000110110011110010110000110000011111001101100100011000100100010010001011001100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out934[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out934, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101011000000111011000101010000010101011101101001110000000010000100001110001000000100101010010011110001111100001000110100100; 
out935 = 128'b11100110011000100000000100000111010110000100000010010110100001011010101001011100010001001001111110010111100101011101110101100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out935[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out935, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011111101110010101000100101001111100001100111000000110000011010011100000110111011000010110011000100001110100010101100111010; 
out936 = 128'b00011111001111110011010100010010110000101110100010011001000001000101110011011111101110100010011111011100010011111011100010100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out936[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out936, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000000001001011100111000010011001001010110101011110000101111100110111111100000011000101001010001000000011000011000001100100; 
out937 = 128'b01010010000101111110001000011011010011011000110111000101101011111010011011011100101100011011001001101010101011011110101100111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out937[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out937, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100100001101111010011110110100000110110100111110101110010110000101010110000100001100110100010001001110001001111000100000010; 
out938 = 128'b00001011110010001010101101101100110000110110111110100101010001011111011010001011111100111010010011110000101001101111110111000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out938[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out938, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100000101010000111111000001101111101111101011111000000111000101111111100111110000100001110011110110110010100111100011000111111; 
out939 = 128'b01111000011110101100110001000100101111101111000000100101001001110010110001011110100110000010110111011100000000011111110010101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out939[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out939, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001110001101010100111100110111000010010110001011001011111000001111011001000000100010011101000100010110110011001010110011010; 
out940 = 128'b00100100011110111011101001101101111011011000001101110110001010010001110110011011000111001100111111111011100111000111001101101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out940[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out940, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101010101001011100101110100001110100010100000110000100001110100000001010000011000110011011110011001010111001011010101101101; 
out941 = 128'b10010101100101101010110001010010011001110101000010101011000000011110001001001011100011000010101011010010001011110001011001111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out941[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out941, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011101110010000110010001101011100100011100010000000010001000011110010010011100010001100010110001010000111110000001011110001; 
out942 = 128'b11100101100001010001101101000110001111101000001110011010111010011001100100011100001100111010000110100011000101111111010101011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out942[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out942, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001011000000111001110001111000000100010010000010001100111111111000101100111011110101001110101110010001110010111000010110110; 
out943 = 128'b00101010110000001101001011001000011010010111111100010100000001010011011111011100101101111010100000101111010101000010011001111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out943[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out943, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100010011110101000101011101100001110101100001000011100101111011000111110011101101111111011010011010101011010010100100101011; 
out944 = 128'b11010000010001000100010101011010110100100100000000110111011010100001110001101101011001001001001100010111100001111101001110110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out944[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out944, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110111111001110100111100011100110100011100000100011000010100110111010110001101101110101101111001001101011110100010011000000; 
out945 = 128'b11111010010101011111100100000000011110001000000100000110011101110001110010111011011100100100010011010101100011010011101111010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out945[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out945, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100011000011000011000011001111001000100001000010010001001000111000100011110100110101010111001001101111010110111100011111101; 
out946 = 128'b01101100101000010101000010111111010010011011101011100111001100111111011010101000111010101011001011111000000011011000010001100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out946[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out946, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010101101111001100110100110101110011001001010111011110101001100111000110110011111100101100101011110111111111010101000011101; 
out947 = 128'b01111111100001101110011001001010001100010011011111111101100101111011110011111001110110100100100111111011000001011100010111000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out947[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out947, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010111000010101111010001110110001111011001100101010010001111100101101111000011100101011000010011111011101100011100101100111; 
out948 = 128'b10011100110010011101011010010101110111111111110011100100101101000110001101111001111111100001111011010001011111000100000000011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out948[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out948, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100110100010000111010100100010010110000011011010111001011111110100011010000001011001100000010011110110011011000010000010001; 
out949 = 128'b11000101100011111010001101001000010001011110010110100000111101101100011100001011011111011111010100010011111100100010011100001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out949[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out949, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001001000100011111001011010111100101011001010110110011010110100000010100111110111100111001001001001101000000011000100101111; 
out950 = 128'b10111100110001100110101010100110101011001100101011011110001000010111001011100100010011010101000101111011100010010111111000101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out950[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out950, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101010001001101010111101111010100110011111001110111000001011000110000101111010111010110100101001000011000001000111010000011110; 
out951 = 128'b10111100011001111110011111011111110001001010010001011011100010001000011110001110011111000011001111011001111101111100111100000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out951[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out951, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001010001000101011111100010000101000100000011010001011101000010111110010101001101100101100011010001111110100010000110011010000; 
out952 = 128'b11001100101100000001000110010111111000001110011101000110010101111001000101001011001100001001111001011111000000110010011010101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out952[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out952, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001010100000101010000100100100111001110001010010111010010001001100110101000111011100000100101000001000010011000010011000010; 
out953 = 128'b10010111100100011110110001001100110001100100000010100000011011011001111011000101010001010000011011100011010010110100000100011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out953[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out953, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011000100110110101010111000011010110100101101110000010011010011111000010110111100001010100100110001001101011110010110010101; 
out954 = 128'b01001111100011011000110011001001001000110011000000100110111001001010010110111110111000001000011101010001011101011111100111101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out954[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out954, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011010010110011100011011101001101001001111001010110010010011001001111101100101110110000010110100111001010001100111100101111; 
out955 = 128'b00011001100000000110110000101111110110100001110000101101000101011111010011011100011110001111011011001001100011011010101110000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out955[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out955, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110000001100111001110101011100100110010111100001000010100011001000101101110000001001100100000100100001111110010011111010010; 
out956 = 128'b01111011001110100111100110000110111110010000110100000111000011000011101000101100000111001100100001001001101001100101100001011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out956[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out956, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000101001101001001010110000011001100001101110000111000101101100101110011000101011100110001100010111011010111110011011011101; 
out957 = 128'b11000011001001001000111100001011010101000011100000111000110011010000011111011110111111111110001010011011111010101010001100100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out957[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out957, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000010110111010011101010001101001011110110111101001110100010010001110001111010110100111011101111100011100110110110110011000; 
out958 = 128'b00010110000010001000010110110101001101010101011000010000000001111001000110010100000111110101100001000101001011110011110000010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out958[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out958, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110101111101101111111100111101011000111111011110110000010100011000101001000100100100011010110111101001111001111001101101001; 
out959 = 128'b11000110101110101011000011001010001100111100001010011101001100100101100101010001110001010100011001000011100101011110110101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out959[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out959, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101010111000111010000011011100111000010101011111110011111001111111011101000001110001001010110111111001110110000111010111001110; 
out960 = 128'b10010101111010001011011001111010000111111011000000110100001101011010100010110000100011110001111010000111100001010001110010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out960[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out960, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111100110001101000110011000111010111010101000000010110100110001011000011001010011010111100000010011010100010100100110101001; 
out961 = 128'b10111101000000100101110000010011000010011001100000110100010101010100101011000010100111101101111000011001010100100111110001111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out961[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out961, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100011100100001111110010010000001001010011110000111010001001011001011111111100110110100111111011000101000000001001000110111; 
out962 = 128'b11101001010110101101111101001011000010000010010000010101100110111110011111011011001100001011010111010100010010010110010100111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out962[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out962, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111101011010001110011110011010001010101101001011111100000111001001100011110101001101010011101010110011100010101111001010101; 
out963 = 128'b11001110010100011011110101001011101011001111111100110011001000110011001011010011101100001000011100010010001110111101111011011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out963[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out963, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010111010101000100101110001001010100111000101001010011010010010111111100110011010000001010001111101101010100011101110001101; 
out964 = 128'b11011010111101100110110100101011010011111000101111010111000101010011111101110101001001000010110011111111111101111110011110111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out964[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out964, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011101101011100111110001011011010010001000011101100110101111011100111101010011110000000011001100001011101001001111101011010; 
out965 = 128'b00110101100000100010011110000001100101100011101111100111110101101000111101101101101100101100100010110111111001011110101001110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out965[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out965, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110011111110100001110011010010011110101100001001100000000111001110111101111001100111000111100011110010100011100101111101000001; 
out966 = 128'b01010100010100000111111110100110010111110110110101110001000111001110011101011011010111011010100011111111110100011010100111110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out966[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out966, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100111011000110001100000110010001100110101111000011100111111001010011110011001110011110110000100101110011011011000101011110; 
out967 = 128'b00010011011000101011000010010110010000010010100101000000000101010010010011010010011010011101000011000110101111010010011100010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out967[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out967, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000010110100001110001100010001000011000000111101010100100101110010010110110111000001110100111100001100011101000100000011000; 
out968 = 128'b10110100011011110001001110010011010100000001011001001110110101000000111101001010111000011101100111010101110000111001000111101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out968[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out968, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001100001111100101000010111101111010000011010000101111001110100101010010101011111010110011100001011101110111111110011100000; 
out969 = 128'b00101011011011100010100111001111110011100100001011001011110001101001111010110110010011101100001000101001010000001001111100011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out969[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out969, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011001101110100110001100100011110011001100001100110100011000110001101110010111101000000100011111001000101101011001010011110001; 
out970 = 128'b00101001100100100111100111000001100011010010011111111001110010000111110010000001010000100001010011110100001101111110101011101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out970[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out970, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100000010111001011110011100011000100101110100101010011001000011111111001010000011101101101110111100111111101010011011111010001; 
out971 = 128'b00010111111111111110010010011000000001111101010110100101001101000110011011001101011101100101100011010001110001101011000111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out971[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out971, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010000001010100101010011001010010011110011000100111110001000000111111101011011000110001010010110101010110100110001010000001; 
out972 = 128'b10110010100101001111100011101101001101010100101110110010011011100000100100001000100100010101100101110110111010111101100000001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out972[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out972, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110110110100100111000110111110010110010001100010001101011001111111001101000100101100100010110011110100100001011010000101001; 
out973 = 128'b10110010010010001101100101001001010001101010101101100110000100010011001100100010100110111011100101011100110110111000111101110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out973[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out973, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110010100100100000100001001101001001101111101111111111000110110111000100000100011010001001111100111000110011111010111110011; 
out974 = 128'b11111001110100010110010111100011000111000000110101111110010101111010100010111011101100111100001010001111011111010010000011011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out974[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out974, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100011001111001001011111000110111101100110101101010101111111001001010111001001100101111010010101100101000101110011111001001110; 
out975 = 128'b11001001010000101101001010101101101011000000111100000110011111111011101001001011111011101101111010101101011100100100111001101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out975[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out975, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011111101100000110011000100001101001110111100001100011001110000000100010101101001011101100110011010001100010010110011100000; 
out976 = 128'b01010000001110010110010100001100010111110111110001110111101011011000100111111011101100111000001000010011100010111101000011001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out976[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out976, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110110000000001011101000000000111111110010010100110010000000011011101110101111110111101111100100001110010000111100100100101; 
out977 = 128'b11001010001011100110000100000011011100000110111011011000001011110101010101111101001111111101110010101100111101000011000000011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out977[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out977, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001011010111100001111011000111111100001111110001010111110010100110011011000101001011000101100010110011001111101111010111100; 
out978 = 128'b00010000011110101000110000000001110011011101100000000000110000010000101011101010110100110011110101001000111111101101101110000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out978[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out978, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100001010000000110000100110100000111110011000000101001101010000010001010110110111000101011111000011100100010111011011110000; 
out979 = 128'b00101010110000000111111011011101101001001011000001100110101011111111100011011000100000110001101011010100001010101000101010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out979[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out979, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111110000100000111000011001000011001101011110111101111000001001010011111111001110010011100001111000110101110111011111101010; 
out980 = 128'b10010001011100011011110000000001010000000000101100000110111111001000000001000101011100100011011011101101111101001111010011010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out980[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out980, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010010111001001101011001101111110001001110010001111000011101110000010011011000010111011010000101101011101011011000011101101110; 
out981 = 128'b10111010000010010111111111011101111101000001000000100101101010110110010001101111000000001110011110111000110001100110000001110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out981[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out981, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101010010010001010100101100011111011000011011100111000011111011001100111010111000100101001100011110100010111011011001111010; 
out982 = 128'b00101101000010100001011110000010100101110100011101100101100010010000000001110110110110110000111001011100011111001110010110111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out982[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out982, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001111001111101011110110011101111011011111000110011011000000111010011101111100011011010010011000001111010100110001000001000; 
out983 = 128'b01000000011101010011011101000100100000111100001011000011001011000011010110101110110010001100010110101110011100000101011110010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out983[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out983, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011110000111011001000100100110111001000011101100101111001101000011100111110000010011011110110111110001001011101010110010011; 
out984 = 128'b11101010010100110010101111010101111010001100000010001000010101000000000110111011001100011001100001011001001010010101110110100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out984[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out984, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100011011010011010101001011011111101111111111111111000010110101110110110111111011100011000111101000101000000110000011111001; 
out985 = 128'b00010000010011000000000110000110010001101010111000101101101100001101000011101000001100101001111111010111000000111010111101110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out985[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out985, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000010101011110010001100010100010000100001110011011011001010010100111000110011000100001011111011110101110011011111100000010; 
out986 = 128'b10111010011000111100001100101110100010100101100011101001110100111011000001111011000111100111010100100001000010001010010000101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out986[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out986, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101100100111010111101111110100100110110110010011001000010110001100110100011011110110011101000001101101110001011100110001011; 
out987 = 128'b11110010001011000001101010110100011111001111000101110100110100010011011111010011100110000100101111011010011111010111100010111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out987[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out987, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110111101110010000110011001011111011111101001110111001110011110010101010111000010000010101110000010001110001101110000111001; 
out988 = 128'b11010001110100111111100110011011011111100100010100110011110111101011110110011001001000110110011100011110011011100010111111101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out988[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out988, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111110101110010011110001110000001001011001011101110010110010101111010111011100100100011000110101100111110000001110000111011; 
out989 = 128'b01101000001011100001100001011001011100101001110000101011011100110011110100000111110000010101011111101001110100110101011100000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out989[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out989, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111000010111101001011000001101101101010000001011001101010010000000110001001101100011100000011000101100001000010010101110000; 
out990 = 128'b00000010010100101111111001011001001110101011101000001101010011100111001010110000110111110011001001110001010010011011111110110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out990[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out990, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011011100100111110100110100001000101100100110000001011101011010001011001111101001110101110100101001001110110101011000101110; 
out991 = 128'b10000010000100000011111101001001000000111110010011000111001100011111000100001010111000001001111110001101100100000010110010111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out991[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out991, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010011110010011011111000101010110101111101001010011111111000000011111100100101100101000011011000110110001001000010111011011; 
out992 = 128'b11101100101100011111100100100100011111000110111100100000000010111010110011101011011000111101100111001101111110100011101011111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out992[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out992, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111100010111100111101010010011100010000000111111010111010011010101100101110100101001001000001011001001101010111000001100011; 
out993 = 128'b00001011011011101111101100001111011000000100011101111010001100011011111010110110111001011010110011000001001001110100101110101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out993[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out993, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010001001000111100011001101011111000001001011101001100000010100000110001100000111010000110001011110011000101011110001011111; 
out994 = 128'b11010101101000111001110001111010100101101110001011010001010010111110110000101010011001001100011100010110001011111000001110001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out994[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out994, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111111100010100101101000010111100100101011001101101101101110000101110011111111110011101111000101000000001111111011100001100; 
out995 = 128'b11010011110000111100110010110011010100000110011110010001001011110010010110111001011110011000010110010110011000011111100100110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out995[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out995, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001110111101101010001000101001100100010110001011101110001101101010101110100000010110111100000001001101111110011111110111100011; 
out996 = 128'b10011110111001010001011100110001011011010010101000000101101101110100001111101001100100011101110001001110100110011011000011110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out996[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out996, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010001110001110110001100010010001000111010100000100000101001110001110011001111001011010110111101111111100011010000000100111; 
out997 = 128'b00101010111110111001101111111001111000001010011110010100011110001111101001101100101111101111000110011110001111100001000101000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out997[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out997, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000110011001111011110101101100110000101110010111000111000011001010101100000000011010000001100110110110000000001010010001100; 
out998 = 128'b11000000010100101001000101000101110011110110110101000011000000110000111001011011001110010111001001101100000110000110010010111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out998[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out998, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101000100011101010111101100000101011001000000010011100010111010111111111011000010110011001000100010101111101111011110011001; 
out999 = 128'b10000100010011010011110111101101001000110100101001101010000110000010010000101110111000111101101101001100000110011011010101010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out999[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out999, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000101110010100110011111000101001111010000010000001101111011110100110110000011101110101010000011100110111001010000101001100000; 
out1000 = 128'b01010000101000011110011001101010111000000111101101101111101010000111011000110000000100100001111011100101000001100011011010100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1000[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1000, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100111010001010011111111111111110111101000010000101011110110011100101111000101110110111011111111010100000011011000001011011; 
out1001 = 128'b11101101110100101110000010111011011100100110111011111000001101001000001001001101011101011101000111111011001011010001010101111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1001[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1001, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000010100011011001000001000110100001111100011101011110001000111100111111010010001101100000011100011110001101101011000000010; 
out1002 = 128'b01000001010111011100100001001100001111101000110110111011110110110100000110010101110101111111001110111110100101001100011001111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1002[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1002, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010011010011000100111001101111010111110010000001111010001000111110111001011010111101111001110111001110001110101011000010100; 
out1003 = 128'b01001000101000110001010100110000111000011110110110010000101001100011010010001101111010101000000011100010000100100011110011001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1003[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1003, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000001011011110001010001100001011011011101001100010111001100101111101101101110010000001111010100000001010110001110001111011; 
out1004 = 128'b00100001011110110010111110111100100110010100111000010001011010101011001111101010011000110010100001110101000011000000100110001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1004[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1004, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011110100001011000110000111111000011001011010001100011001110110001111100111001110000100101011001000110010111001001101000000; 
out1005 = 128'b11100001001001101101011101001001010010000100110110100010100111110001111100110110100101011001100011111100110110000111011000011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1005[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1005, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110101110100100101110100100101000010111011111010111001101100111000001100110000110010111110100101011110111011000110110111001; 
out1006 = 128'b01010001110010010011100010010111101011011011001110110001101010010101110100001000010000010011010011110101111011001011001110110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1006[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1006, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101100011011010110011000111011011110011110111101110010011000011111110110110010011101111101011000101011101001010010110011010; 
out1007 = 128'b00110101011100100010010011101100001001111011110011011110011011001110011111101010000101101011011010010010011001110110010110100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1007[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1007, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110010000001111011001001111100110001110100011110111110000100011001011101001010110110010001101010010011111100111100100011101; 
out1008 = 128'b10100100101101010010100011110111111001010000110100111001000111100010010100000110111101010100100111001110010010011000110011011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1008[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1008, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001010100101010010110010111010111100101000100001010011110110101000101111101000001110000001111001000011001011111110100000101; 
out1009 = 128'b10101010111001001110110000100000100011111101101111001111000101100010001001100010110110000100000001111001001000011011111001111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1009[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1009, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000011000110000001111001000111010000101010000000111111000100110110111101011010110101000101010001100001101010000101010110010; 
out1010 = 128'b10010000010001111110101000001110100010011101001011010001110011010110100000100011100110110010000011000110111011111011001110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1010[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1010, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011001110100000101011100011001100111110110101010100000011001010001110100011010001010011111010101011000001011111001110011101; 
out1011 = 128'b10110110010010010101001010011010110001100010101000100101001011001001111100111111001101011111101101010100111100000000010100001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1011[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1011, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110101100100101011111000110001100100000011010010101001100011000000111100010101110010011111010110000001101010100111100111010; 
out1012 = 128'b11010001101001010011100110111000110110110100110001010001110010101010110011101000111000100101111110001110101101001001011001010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1012[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1012, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001010111110000011000100100010000100011000101111000101011110101001101101001011111110111110111000100001001011111010101010000; 
out1013 = 128'b10001010111000111111000111100000100001101100100010111010011111111100001110111110000111001010111101101111001100100001000100011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1013[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1013, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010011001110111111101100111011110011000110001100010000100010000101001000010000011010000100000010001001011111111001000010001; 
out1014 = 128'b11101110101000011101001000100000111010000011110010000011001001010110011111110111111101000101010000101000001101001100000100110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1014[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1014, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010110110011000011101110101100011010100000111001111000000111010001001001000101010010001011101101011011111101100111101011011011; 
out1015 = 128'b01011111101110000010101110110100111001001010001011001100011001101011010101101100100000010000110010110111110101110111010011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1015[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1015, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011100000100010101111110111100000100101110001001011010101010111111011110101011010010111001001101100011000011011101011101011000; 
out1016 = 128'b00111000111011000111001000111111000101010100010111110000010110110001011001011101000000110110101111011100001011001111111010100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1016[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1016, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001010111010001011011110111100111101011001001110011110101111110111111001001011000110011011110110100100010011110000100101011010; 
out1017 = 128'b01011101010011101111111101011001000000010110010100010100111001101000101011101101011110001101000010100001011011011011011101101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1017[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1017, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011010110100100011011011101110110011111101100001011111110110001010010001101000010100011011111111100110110000001011001000111; 
out1018 = 128'b00001110010111100001111001111111110101111001000000010011000001110101101011100011000000101111001010100011110000011100100001001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1018[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1018, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010101011000000010100001110010000101100100001011011111100000100001011101000111110110010111111011110111101100110110000010001; 
out1019 = 128'b10010111101011101011100010011100000111101101000111011110101111001011111110000001111011011100110011111010110111010001100001010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1019[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1019, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111111010101111110011010100100001100010010011001000010111110111110001011010100110110111100011001101000100111110011001100000; 
out1020 = 128'b00110010101000110110010001110011101101001000011011100110011011101000001100001110011011111010101000110010000111110011111100001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1020[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1020, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001101101111011100100100011100001000100000101000111101001101010111000111000000111000001110110100011101111110001111100000101; 
out1021 = 128'b00111111100001100011110010011111111010111100000011110110001000000000001011011001001011000111001100101000001001110110000010000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1021[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1021, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100111001100101111011010000010111001110000101100100111110000101100110000010100101010111000001111011100010110110100101001101; 
out1022 = 128'b11001100011101011100010111111001101111000110110111110000110110101111110110000011100101000001110100100001001101011100011111100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1022[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1022, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011010110111111111111010101111101100100100110001001011010101101001000101011000000000110100101001011000010101001000001001001; 
out1023 = 128'b11001111010011011100100000011010110111111100100110111110110100100011000000100001001001100000010110000111110110000001111101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1023[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1023, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011100111100010111101010001110000100100001001000100110111011010101111011010011111011001111110011111110100010011100011101100; 
out1024 = 128'b11000111110111011000111110000110000111110011011101011000000000101110111111110011010000011100101001000010010001110000110011011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1024[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1024, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011101011000110111011001110110101000101000111010101101101000001011110101010100010110100111110010011001110110100101010101111; 
out1025 = 128'b11110100101011110010100100110000101101101010100101111111010101110010001111110011101000101101101000101100000001011100111101001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1025[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1025, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110111011111000111111100011001011100011011111101010001101001101101110110111001100000001100110110100100000000000100010001010; 
out1026 = 128'b00011011011010001010101001010100101010010001110101111110010100111011010110010010101010000110101101001100000010010000111000011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1026[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1026, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110011110101100100101100110111001010100100000000100011011101011011010101001101111110111011010010000001000111000010010011011; 
out1027 = 128'b10000100011001101100001000110001001110101001100001010101101011000011110011100110011110100111111000110100010110010111011010111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1027[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1027, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000111011101101010010100111000001110010101110110010001100011110110010001000111011110001010101001100001111100101110000010010; 
out1028 = 128'b01100111010010100111010010010110101110100001100010111011110001010010000011001000010010000101111010110100101111010011000111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1028[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1028, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101111100011110111110000010110001110011110010111111111101011011000111000110111110001011001001101001011111010101101101011000; 
out1029 = 128'b10010100110011000110101101100011111101100111101111010101010000111110010101101011000110001000011000101100001111010111010010011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1029[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1029, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010001001010000011101100100110100001000111111010010011010001000111000100100101101010010111111011111101011101011001101011100; 
out1030 = 128'b01010111110110100101101000010011011001101001100001000100111001110000101100111100110000001101111011101110010110000001100000100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1030[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1030, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110100110001110110000100010001011100011101100010000011111101110000001001011001111100100100101111010000011010010011111110010; 
out1031 = 128'b00001010100000001100011111111111110111101110101011011101010001111000011001110110100010001100101100111011110000011000001011001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1031[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1031, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101101110101110001110111111010011001000010011011001101001010100011001101100111001110101000101001110111110010000111111011011; 
out1032 = 128'b01111110100111011010100111100111010100011111011110010111110001100011111111101011001111010000110100010010110010111111101110001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1032[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1032, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101101100111001010100110101100010110101001110000111110011010111100110011011100011000100000010000101110011000001101111011110001; 
out1033 = 128'b11000001110000111011001010010111110000111101110010100111011011100000101011001100110111110100010100001010100000111011001100100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1033[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1033, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110000011000010001001111101110101000101101000000001110100110000011000110010101000000010100000101100110000111010110101001001010; 
out1034 = 128'b00001110101011011000100010101001101000101100001000101001010100111011001010100011010101000110010000110000011001001001101101010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1034[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1034, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100000100000001111001000000110101010000000001101000000011100111111101110101110010110101100100010111010010010111111010100100; 
out1035 = 128'b10011100000010100101000001111001111111010110000011010111110001100010010110001100001111000001011011101100100111001101111101010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1035[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1035, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000011110111110010101000100001100001100001001110111101100000001001010000011000110011101101111101011100011100011001001110110011; 
out1036 = 128'b00100100100011001101001110111011111001101101110011111111111111001011001111000100100110110111110011111011011010000100000010111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1036[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1036, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111001000011010111011010111011010001001111111110011111001101100010110001100110101101001010011000000010111011011010111011111; 
out1037 = 128'b01011110010111101101010000111011000100100010010100111101011000100111000100010111010001100000101110111110110010011110011101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1037[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1037, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000010001101100100001101000110111011010010010011001110010110001011001010111110000111100110000111000001000100010001000111010; 
out1038 = 128'b10000000101110100110101010011101110110010101001000010111000001000011010111110010100101010111001111100101001001000110101110001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1038[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1038, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101001110111011001110011000101100010111001000011011011110101101000101010000111100110100001010000010110010100011000101100110; 
out1039 = 128'b01010000010001100010000111111001100101100000111100100110001100000010101011010101001000100101100111011010100010000110100001111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1039[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1039, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100110011011010110000011111000100011011110001010011011110011110001110100011100110001100000101110101000000010000111111000011; 
out1040 = 128'b00100001111101101010111010001100100010010100101000101011011010101010000100011101111111001111001110110100010010100101011011010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1040[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1040, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110101101101010011101011001001001111110001100000011001010011111110111010110000110111011000001010100011010111100000100110100; 
out1041 = 128'b00010110100000111010011111101111010110111001100100000111110010001000101100110001001001111100100001110000010100001110000111111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1041[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1041, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000010110101101111001100010100111100000110010110101001000000100111001100101000001100111101101000001101010110001111001101110; 
out1042 = 128'b00101001110100100001110001110100011111001100111011011000000010000000011101111011111000101011000110000011101001000010010101010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1042[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1042, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000000100101010010101101001101101100011111111110111011010101000111111001100110101100100110110111100101001010000100101101010; 
out1043 = 128'b10001101001111010010011100001111111101011100010101010001101001010111110011101111010000100011110000111111100010011101000001000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1043[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1043, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001100001001110010011101011011001011101110001000100111111001011111101101100010111111100110100010111111000101010000101010110010; 
out1044 = 128'b11101111111000010001101110110111010100010111100011011010111110110000001101000101010100101001110101010011100001101100100101111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1044[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1044, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110100101000010100111111010101010100100100101100110011101110010010101001001101101001001111001001101110001010100010100010100; 
out1045 = 128'b00010001100010010111110011101001011000101000000101010101001010000110011011001010000001111111001000110111000010010101000001011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1045[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1045, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001101110101101001000101000110000101010100001011111100111111100000111000010111110000110110110101110000110011001010000111111; 
out1046 = 128'b00010011011010111000010101111001011011101011010101101001110011000101010011011011111001000010110001010110110100100011011100101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1046[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1046, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000011101010100101111010011010010011101001000101100101110000100100010011100101010100110111110010000000001000000001001010011; 
out1047 = 128'b11101100111110101111100111111010110011010100010000010111110111110101101001010100111000101110000000101110011110001111110111010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1047[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1047, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001010000101011100100101101000100101100001111001001101000110100111010100100110010011110101100110110000011110001110101100001; 
out1048 = 128'b11001001110101100110000010010110111101000000011011011011100011010011110100001110111001001010111011011111001111010110011110000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1048[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1048, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101111111100101100001100011100001011110011111101111111110000000011000000110101111011001111111011100000000111110101111100111; 
out1049 = 128'b10110110111100011000000001111001110100000100001000100010101100000111100001000011111010110001110001111111100101010011010100101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1049[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1049, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100100010110001100011111010010101100101100110010010010100000001111001011011000101101101000010100010000000100011110001001110; 
out1050 = 128'b10010100000001111010110110101100011111001101100010100100000011100110001010110100100110101101100100101000111110001110101101100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1050[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1050, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111001000101100011111111011000011110110101010011000011001000001111011011001100001111110011110011101010110101011100010001001; 
out1051 = 128'b11001100001001000000110101010001110110100110100111000010011110011001011010101101111100010001011110000000001000000000001101000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1051[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1051, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011000001010100101011001101101110110110101000110000101110100011001000010111100110100010101100110100000100001111000000000110; 
out1052 = 128'b00000100011100001100111001110010111110111100001011100110000010101011010011111000111000011011000101100011100001000011001000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1052[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1052, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110010111001011010100111110001011011000111101101011010101011100111000001101011101000011001110010000111011001001011110110010; 
out1053 = 128'b11100110001101010110111011001101010000111101111111111101010000000110111000100011000011000110100110110101110100001101101111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1053[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1053, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100001100010100111010000100010010000110101101110100011000010110011010000100100100010100100101100111111010111011110000011101; 
out1054 = 128'b00111001001010001111101110010010111101010110101001111110110110011000000101000101101010110110000101011001110010110111000110011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1054[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1054, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110011100000010111110011101101100110101011010000011001000111010101100100111100000110101111100010001011010001011110000001111; 
out1055 = 128'b11111110110111101001100100111101000100101101100101101000011101101110110000011111110000100001111011101101001000100001100011011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1055[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1055, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000011111110000001111111010011111001110111100110111100010110111011001100001110011111101010001111100001111010111110000010100110; 
out1056 = 128'b10010000010101011111101000101111000011100110010111010001111110100110010001100111100001100100000100001000000101000011000011101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1056[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1056, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101011100010110010101101010011010110010110111100000001001101100010110110011101011010000010010000101001111001111010001100000; 
out1057 = 128'b10101000000010111010101010001000100001010000010010111011010010101101100001100010011100110001011011101100010010100010101000110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1057[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1057, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001010111110110110011100110110110010100010110101001100001011111110111010001011010011110000011111000001000010000001111000010000; 
out1058 = 128'b11010011011110000100000100011000001100110010110000001001111111010110111110110100111001111010110111000110100011111110110100001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1058[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1058, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101111100110101110001111100000001101101001100111101111001000110001111011110111100111001000001111111101010111110100000101110; 
out1059 = 128'b11001000011110010101111100101110000110001001010101111000000001000011000101010001100010111100111010000000100100001010100010111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1059[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1059, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111001000001101100011000001111000001111101110010001001011100101101000101010001010010011111011101001101001111010011110011000; 
out1060 = 128'b01110101110010100001110010001111100101000010110110110101110000010110100000001111000000011101011000001110101111011110000001011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1060[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1060, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101011000110111001010110111110111101101011110110010110000010010011111001101010111011011110110101001110001100100000000111010; 
out1061 = 128'b11101101010110111011111000100111110110110000000011110000100110101010101100011100110100111010001111001010100000010011111000111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1061[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1061, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101010100100100011001100000111001101000011110100100001011010010111001001110010101110100000000011011001100000111010100011010; 
out1062 = 128'b11000110101101000000111011100100010101110010000001100011010111010111100100101100111111101111101101010100111101100111111000100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1062[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1062, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111110111111110010010111111010000001111001101000100000010101111010010101101100000110110001001110101011001100010001100101110; 
out1063 = 128'b11000101101000010011101100100011111110101010110000000010001001111101110111110001001100001000000010001011110111110111111111110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1063[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1063, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001111011110011001110101111110000111110110101101011101111000110000010111011110011110101001011001111101111010110001111010011; 
out1064 = 128'b11110010111011111000101110101100000000011101101100000011110101111010010101010111001001001101011000111010110111000100011111101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1064[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1064, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101100001111110110001011011010110010010110010100111001110010011111110000101111011000010111111001101001001100100001010111000; 
out1065 = 128'b10100110000010111111000110000110111101101101010110100000000001011001000111101000111101110101010001001000001000110101110001110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1065[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1065, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010000101100011111011111000101100101110101101001010000000010000111001010001110111011001101011111111000001010010010111010001; 
out1066 = 128'b11101010001000000100110011010100100100110000001010101001110100100011010011001001110011110001010001011100101100001101000010110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1066[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1066, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001001111000010010101011101110001001001100011001101100011001110000100001000110011000100011100011011000001011001001011110111; 
out1067 = 128'b10001001110011000011000101001101111100101000011111111011010010010110100011111001000101000000100011101111100011011000000001110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1067[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1067, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101010110010000100110111000001101010111111011111011011100100001011011111001110011000101001111010000110110000001110000010000; 
out1068 = 128'b10100100010001101111111111111011111100101000101110100011111110101100110001011100101010000001010011101111010111111111101110010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1068[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1068, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111001011111011011111010100101110101010000100010101101100010111101100011111110010010011001111110001101110011010100111111010; 
out1069 = 128'b11100101111110110000011100111110001110000001111111000000111111100111011110001011100111010010001011111000110100000010111010001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1069[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1069, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100010000110111010011000110101001001101001011101110000010011110101100110110100111011011000101000011101010110101110110000011; 
out1070 = 128'b11010110010100110001011000101111010000111000000110011100000001000011110111100010010000001001100111110011100001001101110101000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1070[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1070, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101001001000011100101100100101100000000110010000010011010110101110000011110010101001110101101111010011111001110001000000111; 
out1071 = 128'b01110101111110100001001001101011110110000100011101000010010111010111010000110111011001011011010001000100101001000110000011001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1071[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1071, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001000011100110001110111010010100010110000001001100100100000110100111010110001111110111100101001010100101110101001010101000101; 
out1072 = 128'b01010001110110010000010001110011111100111011101100111111100111111111010101111110001100111000110100111110000101011001001000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1072[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1072, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000111100100110000010111101000100010100000010101111111110010011011100001111001100110000010100101011110011110111011001011001; 
out1073 = 128'b01001100010011101010111001111000011000111111001100001111110111110100001010111100101010100000110010111011011001010100010001011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1073[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1073, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100000110110010101011100010101101011101111011011110100001001010011000111110000111011011110110111001011100101100010011101100; 
out1074 = 128'b01101001110001100011111000001101011111110010011110000101110110101000111011101001001101110100000010000011111011110111111100000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1074[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1074, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011111101001001000111011010111001101000010111111011010010111101011110111101110010010000111111110100100110001010001111101011011; 
out1075 = 128'b01101000001000000101011000111100000000100100010010001000010001101110111110101011010101110100010000000111101101100110011010100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1075[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1075, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110000001111001001101100101100110110101000010111110011000100110111111000101001111101100001001100010110111110010011101010101; 
out1076 = 128'b00010001101111100010110000001111100010001011101110101110100101111011000010010010001000110100110110001000001110011111101000100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1076[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1076, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110111000110001100000111011010000100010010100101010110000101000101111001011100110000100001000100100101001111010100110001100; 
out1077 = 128'b10001010111101000101001100010101000101010100001110010011011110100010100110011100001110101010111101111100011111101010010110111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1077[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1077, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001000100001001100101100000100000001111010111110100001011000111111100010101111000110011101110101111110110111010000000001100; 
out1078 = 128'b01011100111011001100100010100111101110001110100000100001000100101111010101011001110110010101001010111101110111111000100000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1078[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1078, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001110001110011010101000011010100010001001111100101100000011100001011100100000010101010001111001011100001110010111111011001; 
out1079 = 128'b11010010111001000101100001101011100000101000101110000010000101111100100010101101011100000000100011101000000011010110010000010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1079[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1079, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100001010100010001111001001010000110111010110011001001011011011110010111100000101001111011101000000111010010101011000110011; 
out1080 = 128'b00010111001001100000101001010100101010011101100011101110100010010011001000010001001100000111100011110101101011000100001110010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1080[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1080, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111101101100101010101011100101111111000101110101000101011101101001101100000000111000111111000001011011010101111101011101100111; 
out1081 = 128'b00100111011000001011100010001011000000100011010001010011101110010110101001101011001000001110101110100110111111101011001001111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1081[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1081, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111011001010110011110110101011000100100010010110110001010011111110101101111010000011001100110101001001100110111010111111101; 
out1082 = 128'b10100000111100100010100101000011111111110101101101011001001111001100100101001101001111101001010100010100001111100011101001011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1082[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1082, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100101100110111011000101111101111011011001100011100100011111010011010001011101111101001001011100110100000111110100110101010; 
out1083 = 128'b00000110101011010001101111010001111000110100010101011010111011110010111110000010001001011001010111101010001101011000101010001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1083[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1083, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011101011111000010111100010011000110111110101000110110011010010000111001011000011101000001001011101110111111001010010000100; 
out1084 = 128'b10010111010101010110100101000001111110101110111111111011011111100010101111111000101001000000110001100010001010010000000100100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1084[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1084, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111001111010110110110101000111011110010100001100110111111101100011110101100011011011011011101110010101001111011111111001100; 
out1085 = 128'b01111011001010000000000111000010000111010011100111111011100110000011100101101011001011001001001000001110110010111101011000111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1085[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1085, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011110011001000000101100010000100010100010111110000101000110101010110001110110000010010001100101010011110101110010011011100; 
out1086 = 128'b11100100100101001101010100110101100100111100000000000010000100000010001101000101011010000111100001100000101110011001101010110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1086[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1086, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001010011111010101111101010001101101011111010001011111000101101011011000111000001100000011011101001111010001111101110010010; 
out1087 = 128'b11100000000010001111000100011001010000111101001011010000110011110001101001100110100010100101010101111111100010011000011000100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1087[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1087, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011111011010001000111111010110101101100000101011010111101001101001010111110010111001110010110101111110011101101111010101010011; 
out1088 = 128'b00001001001111101111111110000101010011011001100011000011100000001101010100100011000001110010101011100100000001010010110010000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1088[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1088, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111111101001100001100101001101001101010101100111001010100101010010000001011001101000011101011100000001101110000110010110110; 
out1089 = 128'b01000010111001111011011001011110111100101111101010100000011010100011000000101001100111011001100001100011111001110011001101111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1089[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1089, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011001101101010010111100110110101111111101001011101001000101100100110111111101101010100110000010111110011011010001110000001; 
out1090 = 128'b10111011011000110100100010001101010110010001001110100101110111111011010010000100001101010100111100001101101100001010000000001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1090[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1090, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101110110101111110001001011010110011101101010001000010010011100111111111101111001111010000011101100101001111000000110011001; 
out1091 = 128'b11100010000011011101001010111000100011110010001000001100011000011000011111101111000011100111111101001010001001101100110010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1091[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1091, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100111100001101100010011100100101100100110001001110000011100100110101010001110110101111010101010001100101001011100001111001; 
out1092 = 128'b10111110010011011111100111001100011010110010010100111101001100000010101011001101111101110101110101001010010100001001100011100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1092[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1092, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011101000111000011101101011110111000001110011011110111001001111000011110010111100000101000001100100001111100000011111011001000; 
out1093 = 128'b01011000100110000110000000110011101010011011101101000110010001111010111111110000101110111000000001111100000100101100111010100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1093[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1093, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010011010011011000011010101111000110010000011001100001101000000111010001111000111100001010010101000001001001100101011010111; 
out1094 = 128'b00111001001111011001001001111111111000000101100011010100100011100001011111000001101000011000101100111001111011100010011111010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1094[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1094, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101010011101011101011010101001100110101011011110110111111100100010101010011100101101001001011011101000010111110110100001001; 
out1095 = 128'b11001001001100001011010101100100101100011011101001011100010000110010001010001111111111100110110011010010001010011100110111100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1095[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1095, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011110001110100100011110100011111101100010011111011111000111110010001010000111111101000010110100101011010101111101001000001; 
out1096 = 128'b01101110101111100110011011101001110100001000101010011101100010100100001011111110101101101111110111001000000110011100010010000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1096[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1096, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101110011110000000110010110011000000000001110110110101100101110001011001101101011101001111101101011101010000111001100100100; 
out1097 = 128'b10010100101111111111000110011101000000001111001010011100010111100100010001000011101010001110110000100001000000101100100011101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1097[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1097, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011011001111100111101100001010111000000000011001111110001011000110111000100100110011001001010010111111110110111010101101011; 
out1098 = 128'b11100110111100110010010010111001111111101001111110011010011010010011001010111110111010101000101001110000010110110001011110101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1098[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1098, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111100111001000111010100111011001101110010111011101101001110010011100110100001001111010111101100111001110001000010100001000; 
out1099 = 128'b11101000111001010101001101111001001100011101111001111110101100010101100111111000001000100101010110001100010111010100100001110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1099[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1099, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110000101000110010010001001000100100010100000111101000111111101010100000100011010001100110111110111100101001000011000000010; 
out1100 = 128'b11011011111011011110100100011011101001100110111010111100011001110000110001001010001101010100110011011001001110010111111111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1100[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1100, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110011100100110001101001011111101110111111111000010001111111000011001100111111111101100010011011001101110010100110111010110110; 
out1101 = 128'b11011100011010111101101110101101110011010000001101011000011000100111001100000101010101001110110100001110001110100000010010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1101[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1101, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001010110000010101111111111010110101001000011000100111101101101001011110011100010011100001100011010101111110100011100000110; 
out1102 = 128'b01001010011011111001111010001100111111001011000100110001110011001110000100001000101100001011000010011011000111111011110100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1102[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1102, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000011101110011010010001001110111000001000010010101011101000110110110100100011001110101101001001110011011100010010100110010; 
out1103 = 128'b11010010100001011110101111110100100011010010101010100001010101111100000011000011111000011110001101011010011011010000111101011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1103[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1103, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010010001001001100101100110000000101000101001111101100101011111110111011111001000110000101111110000000111110100101100010100; 
out1104 = 128'b10000001100000001011100011100101001101111000101010001101100010010101001100101010101110111000011011000010101010100111011100110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1104[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1104, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100011010100111101101101111011100110111100101110001011000100111100100001000111000101010000011110101110001111111110001110111; 
out1105 = 128'b11001010111100110110001011101111101100110111011110000001101100001111101110110111110001001000011110111110010100001001110011011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1105[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1105, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101110101100010001001001010101010111001001011100111100111101011110000101101100100100010000110110100011001001000101010011100; 
out1106 = 128'b11111110011100101011100010100001010111100001000010000010101010001111101100110100101111000100010000100101111111010110100111100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1106[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1106, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101111111001110010100110010010111100001101011101101101001010010101110110101100111101100010000001010101010111101110111100000; 
out1107 = 128'b01010010000010110100000101111010000101111011111011100011001010101110000110110010010100010100110110001110100100100111000111010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1107[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1107, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011111111100011011010011010111100000100011010011000100000011111111111100000001111110000000100100010101010001110000010011100; 
out1108 = 128'b11111101101001011001011001011010000011111110101111010110101000101000001110001001101111000111111000111010011011010101111101010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1108[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1108, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001000110011001010000000100011111001011111001011000001010101001101110011100101111100010011101000100011100000100110101110010; 
out1109 = 128'b00100110110101010010000111010101011000011011111100100000111001100001111100010101000001010000010011100110110110010001101110001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1109[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1109, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100010010001100011011011101111010000011100110001011010001111110011100110010100011100110000001010111010011100100101011100001; 
out1110 = 128'b00110001100000001100111101100101010000111111011011110010011001111101011010000011000101011001101110000010010010110001010000001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1110[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1110, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100000101001100101111101001000100001000011001101000001101000101000001100110110101000110001011111101001110100111011101000111; 
out1111 = 128'b00011001111001111110001110101101010001010110011001101001011000100011100001100001011001000111101100100100010000111001001110111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1111[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1111, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100101101110110001101101100111101100111011000111111100110011111010000011000111001100011110011010000000101101101111000010101; 
out1112 = 128'b10011110110101110110100000111000000011110010111010111010111011111111111100011110010000101010010110111101100101001000101011001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1112[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1112, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000011101011000100000111010010000111110000100000101100001000111001101001001100000000111111011110001101100001101101111110111; 
out1113 = 128'b00010111111110100110001101101100100001101111100100101010001001000000001000011110011000000100100101010010111000010010100010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1113[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1113, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100110001011010111000010010110101100111100011110001011000010011010101110111001001101110111111101100011111111110000100010110; 
out1114 = 128'b11000010100001010110110100000111001001100001101010001110111001101101111101001010110011001011001100001010110111101100001001010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1114[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1114, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101011010111101010001001100001011111010111100100000101010111010001100000001001010010000010111001100110001010101111101110101; 
out1115 = 128'b00111100110001001000000001110101110100000110011110100110110000110100101101010100110111011010000011111000110010000101110001001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1115[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1115, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001111110000111001001010111011101010101000111011111010100100100001100011001000101101110101110101100001001010010011000010011; 
out1116 = 128'b00100111010111111110010100000111010101001001100111011101010001010010011101111001110001101100010010110000110100111110011000000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1116[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1116, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110011111101110010101110100110010110011111011010111010000011111001001101110010111001011110010110010011100110010011100011110000; 
out1117 = 128'b11000000011110111111101111010000100101100100100011111100010000001010001101111111010010101001001111000101010011010101100011000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1117[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1117, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111000101110101101111000101111011110000111000001001011010011110000111100000110101000100101101010011100010011001101001010110; 
out1118 = 128'b10010100000010000001100010001111110101011010011011001100111000001111010011111111111001001010011111000000100101011001011010100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1118[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1118, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110111011001101001001011101100001000001110101001001110010101100100000010101110110001110001111100000101101100001111000010100; 
out1119 = 128'b10000010111001001110001110101100010000010000001110010011001100110110010000111011111001111001011011001110001010001100100010111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1119[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1119, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001110010100010100010001001101111100011001000001101101001000100111000001110100000000000001010111100001011001011110010101000; 
out1120 = 128'b00001011110110010000111001101001111110111100100010011101111010011110010110011011011011110101101100101011000000111010011100000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1120[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1120, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010100010100011111010001111101110010111101001000111110010010001011001110001011110001000110010111111000111101001100010101010; 
out1121 = 128'b10101111001011000011110111010011101011110110110100011001110110000111111100100100011001010101000001100110101101111000010010110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1121[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1121, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001001101001110111111110100001101101101010100001110000111101100100010010000001010110010011111011101001001010101111011110010; 
out1122 = 128'b10000101110110011000010101000111001101100111010110111001110100001011100111001100000000000010111111101000010100110101010011010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1122[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1122, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011111000110101110100101000000010101010011101001000101110100011000000100110110000010111110011011001100000010100010101100101; 
out1123 = 128'b10100111111000110001011111011110011011000100001001011000010011110100111100100011111000101000100100011111110100111010111101101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1123[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1123, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001001010001100111100101100111110001100101011001000010001101000100101110101101110010101001101011001110010001111010001111010111; 
out1124 = 128'b10110010001110000000000101111111100001000001000000000100100001010001010010101100101110001110010001000101110100111010010111011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1124[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1124, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110101001000100110111111100111101110101100100010110000110111011011001100110000100010010001101101100101001100100111101000101; 
out1125 = 128'b00110110010100001101101101100111001100000101011001011011010101000100110010111011101100101010000110010010110111100111010110010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1125[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1125, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101011110111000010101011100100101101101101100111110100000110010011000111101011001110000111101111001110010010001001110101011111; 
out1126 = 128'b00110001100101101101000010011101110101110000001110110110011110110000101000001000101010100011011101001111110110100101000011100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1126[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1126, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100110111000010100010011100001000100101101111101000100001101101111001111001010001011001010101100101011000101010100101010111; 
out1127 = 128'b10010010001011000111000100010110000110011110100011010101011010000111100011110100100111000100111101111000101000001011011100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1127[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1127, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101010101000101011101010011001101010011100110010111001110110000111011101101000001010001111010000011010001101100100111001111; 
out1128 = 128'b00001011101111010010111110000000100000000110100011100001010000011011101010110100111110100010101111110111010100001100010101100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1128[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1128, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110111000010011111111111001100000110010010101110110111101011010100010010001111110110001010110110110001000110100000011110001; 
out1129 = 128'b11111110101100111111111111100000000101011111001010000110110111101001101111000100111000101110100101110000110100100000011111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1129[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1129, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001111110011100111010001110010010110111000111010010101101011011100111110010000111101000110100000110001110101100110111111011; 
out1130 = 128'b10111100100001100011101011011001010110101100101000111100100111010100101110100101110110011001100011000011111110001111000000010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1130[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1130, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110101111010000110101110000000011101110111010101001001010000111111110111111100111010100011101001100010000101001101110011000; 
out1131 = 128'b11111000100110000010101101100001001110100010110100011100101101010101010110101101101010110000111000001101000010000110110001010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1131[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1131, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001100100111010001010100110010001001011100100111011100110110001010010010100110110111011010011010010101010001110010110000111000; 
out1132 = 128'b00101011001101101100110100100011111111000001110100000110001111110001001110101100010111001001010100110000100000010001011110011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1132[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1132, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101010010110111010011111101011000101100100000010001110100011010101100000000110110101001010000110101010000101000001110000110; 
out1133 = 128'b11100011011111011100101111001001001000010011101101011010101000001110100100101001001001101101010100011011110000001101000101001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1133[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1133, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110000000101000100101101100111010000101100101001101011111001111111101111110101001010000001001010001111110000011101010011100; 
out1134 = 128'b00111010100110000111010010100000100001111001001111000010100100011010110011110100111101101011010000101001101000010001110001110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1134[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1134, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101110110010001100101100010111000011101110011010101101110111101101101111001101101111101010110000101100111110101001101101110; 
out1135 = 128'b11000001110110001001110011100100010101011101001101111010100101010111011011011111001001101101110011010110010010001101011110111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1135[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1135, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101101010000101011001011100010110111110100100100001011101100111101100100000011101001010010000101100111010101001010110100100; 
out1136 = 128'b11010001000001010001011101101110001001011011001011001111110100001100111000110010100101011001110010000011101110011111110000010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1136[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1136, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001011100010010101011010011101101111010110001100011000110010000011011101101001111111001011000010000011000110000100010000101; 
out1137 = 128'b10001001111111100000011011101000001101010000001001000100001100001011011101000101011101001110111010011100110000000011000100010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1137[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1137, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101100101011110010111110000010111001001010000001101100010110011001111010010110000010001010011011001001001100110101111000010; 
out1138 = 128'b01011100010111110010000110101000111010000111100001011110111100000110001011110000010000000011100110100101110011011011001101110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1138[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1138, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100101100111010001111110100010010101101001111100001011111011000001100001011001110111100011000101110100100101000001010001101; 
out1139 = 128'b11101010111101100011011011100001101010110111111101001101101011110110000000100101111011100011111001011111101110000010111100000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1139[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1139, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111101000100110001000100001001110000001001101011101100110101000111000101010101001111011110011010011111011011100100101000001111; 
out1140 = 128'b10010011000011011010010111000101101111000011000001011010001100111101011011010100000001001100000011101000100001111111001100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1140[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1140, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111100011010010010010100000010000000110101101101101011111110101011010001011010111000101101001000001110010001101111001111000; 
out1141 = 128'b11001011101001011011001101110111110011100110110101101000000110011010011101100000011000111000010100100000001010000101001100001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1141[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1141, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101010110110010010111100001001010000010000000011100101101000111101100000010000000010100101000011011001000000010110110100101; 
out1142 = 128'b00010001110110100000111000111110010101100011011111011101001010111011101010100110110011011101001101011110101100100011011001100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1142[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1142, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011010001101111111110011010000011010100000110010110000011001011001101110000100101100011101001110110110111001100011011110101100; 
out1143 = 128'b00101011011111101110110110001000100010001101100110111001011110111001001001001101010010001111000010111000000000000001111101000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1143[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1143, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000000001001001111010000110010111111100000010101010001010010001101100011111100000001001010000111010000011010010010010110000; 
out1144 = 128'b10100100100100100111001001101100000010000110100110001011011110001001110001011101111111000001100110100100110010111000100111000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1144[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1144, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000101111100110101011100000111111010001001111111000111111100111001101010001011100100100000001001100000000110111010110011100; 
out1145 = 128'b01101000011100100000001100101000000100000011100101011101100010001111101101100111001111100000011111000110001010010101101011001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1145[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1145, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010110111010101000101000010111000011110001010010000001011100001111000010100000110001011101111011101110011100000010010001100011; 
out1146 = 128'b00001010001101100100110111000001110100100010010111010101110011010011110100001000011001010001000010000011101111111111101100010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1146[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1146, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100000111001011110110100001101011000000010110011111101111011100110010111100000101000011111100010100010001100101011011001000; 
out1147 = 128'b01000100000000000100100000100110010010101110011101010001111100101110001100000000000001011010110110001110110101011101001100101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1147[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1147, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101010001111001010011100010010101101011001111101011110001000111101011000111111000100000010000001000100111100101100100011001; 
out1148 = 128'b00001101001111111100001111111010001110010001010000111001111100010100000111100111010010100111101111010100011001111000101110111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1148[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1148, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101010000010001100110011110100010011001000100010110010011100001110000000010100011110100100101000110100001001101011101110000101; 
out1149 = 128'b00101111100111011011101111001000011011100111010001111001110000001011100111010111100011000010111011110101100010110101000100011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1149[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1149, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001001110110111000100101100011001110000010001011110001111111000111110110001111111001100111110010010100111010101101110110001; 
out1150 = 128'b01011101001111101110111101011100111110101001000101100001001111010111010000001111010110111110111110001011010101010100100110100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1150[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1150, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111110100010101000110010010011001010111111010111010011001110001000000011010100000101000011110011011100100010000000000111001101; 
out1151 = 128'b01101111101110101011111001001101000111100101010100001100101011001010111011001001000101010100101001100010111001101000100100100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1151[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1151, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101100110001101100000011011110011101000100110000111101101010101110110001001111100011001110011101111101111111011101100100110; 
out1152 = 128'b00100001001010000111010001110001111000100100110001011000011111111011101110001111100111000010100001110010011111100000101011110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1152[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1152, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110101110011011001011001010000010101101111100000001111011110001010100011101001101000111011000001101111001101111101001101001; 
out1153 = 128'b11010001100011001000110101001111101101011100100001000000000000100101100001100110100011000011001101010110101110001101101111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1153[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1153, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111001100011101101111010001010000100011111111011101000011100110010000001101100010110101010101001000110000011000111010111000; 
out1154 = 128'b11011010011010011110010000111000110011001001111100100011101111010010001010001010000011011010011100111011100101110010100011110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1154[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1154, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100111010110110000011110011010111001100111110001001110000011011111111101111100100111010110111101001011111010010110100110001; 
out1155 = 128'b00000110001011010000000000000100001010110011101010100011110010110100000110001111010101101111010100000000100101101111111011011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1155[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1155, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110100001110100000010010111111001110111000001110100100111110000011011001100101000010001000100001011001101101100100101001011; 
out1156 = 128'b10011100111010101110011110000000001111100111011110011110111001000001001110100110101010000001001010100001011011000010010100110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1156[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1156, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101001010011100110101011100010101110010111011000100110100011111111001111100001100110001000101011110110100010001111001000001; 
out1157 = 128'b11111000101100110111100000111011010100010000101001101111011100111001101010011001000100000110101011111100010101110000111100011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1157[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1157, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011001000010001110001111001010101100000100100100100001111011100101000001010111010000110010111011001011011111001000110111001; 
out1158 = 128'b10101001110111010100001000001110010000000101010111001011111100011010101100111111100111011100101101011100101011010000010001110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1158[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1158, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100111000000000010011101100011011000110111011101101110110000110100100111111010110111011110000011100011101101000101111011010; 
out1159 = 128'b11010000101000001111011101111010000101111110000100011011001100110000100000000111111100100100101110010011111011011000000100011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1159[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1159, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110001001010111101111101101100111110110101111111000011110110011100001110101100011110011000100000000101101001101101001001100; 
out1160 = 128'b01110101111010100011101101100010011111011100011010101000111011111010001000110111000001001011100000011111100101001110000111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1160[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1160, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001100011100101110111110110101101111010100100010100101001111111110100110011100001000010100101111001000011101000001101001100; 
out1161 = 128'b01111100111111011000100011010010011100011001000111111010000111001001000101100000101111010101101110101010011101011100010111111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1161[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1161, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001101111111011011001000001111100011001010011001101110110011011101011100000111011000100100000100100101001001100110100110010110; 
out1162 = 128'b10010111011001010011100100010110000100100000010000010011110111011011100011011010111110011100011110101101011110001001010010011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1162[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1162, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100110100111001110110010011000101001010111010110101010110010110111100001001000110100100001101110110001010000010101000010101; 
out1163 = 128'b00101001001000000111010100100111100000110101101110000000010101100100001100011110101101111100101001000001101011001101110100100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1163[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1163, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111110110001001101100001000101010100110000101010010100100000101010100111001000011101001101011011111001001011000100101010110; 
out1164 = 128'b11110101000000010110000000010110001110101000001000011010101110110011011100111001110011111100000110111111001010110100110011111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1164[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1164, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011010011010011001001101000110000100011001011010000110001010100100110010000010010110110010010001010110110011110110011010000; 
out1165 = 128'b00101011000000011000000010111110001010111000110110111111001000100000100111101110110101111110110010000011011101010110010100011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1165[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1165, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010011011100110111101101111000001011010100111001111011011101001001111010110111010011111111001010000110001111100110110001001; 
out1166 = 128'b01110010000010000010111100101111000001001000010100011101010011111101100011010101111010000110111001110100110111010000010110100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1166[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1166, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111010000011000000111111101000101011100110001011110111111011000101110111000100111010010001000001010110111001011100011101110; 
out1167 = 128'b10011111111100100011100100011000101110100001110110110100110110100110010010101001111101101011001000100100010011100110100000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1167[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1167, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011110101010111100111011110001010010101011101110010101111010100001010001110001001011011000011101000111100010001000000110100; 
out1168 = 128'b11011010011011111001111111100000110001101010111010011001001001011110110000101011100001011001001111000000010111010101010111010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1168[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1168, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010101101000111010010011001111000011110010110001110101101100000101001001011001011101100100111011111100011011101001010000011; 
out1169 = 128'b00111010000101001101101111111010111100011001010001001010011110101000111001111000101100000100110011000000010010101001100101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1169[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1169, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000000010000100110101001101100010110011011010101000111100011000101110001101111001111101011111010110000000011101101001001110; 
out1170 = 128'b00100101011100111000101111001011000101100110101000001011010111101010110110010001111110000110010001010011010001101000001000100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1170[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1170, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101001011100010100110100110010010010001010110011111001101001000000110001001110110101011011110000011001100010100111101111010; 
out1171 = 128'b10101011001000111101111000100111000000110101011001111110101100110101000000001001000100110000000011011001011100111111010001100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1171[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1171, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010011101000011101111001110010000101011011110000010100001010011010100101011110101000010101011011110100110111101001111100011; 
out1172 = 128'b00000100010000001100110100010101111001111111111011100000101010011110010111101010010010110101100011011101001110100001001000001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1172[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1172, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011101100010011101011010110001011010100010110101000011010001100010001011100101000101010111110100101010101001100000101110011110; 
out1173 = 128'b01000010111001000001101000000010101010100100110111011101011011111000010000100111010001111010011111000111000010110100110000101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1173[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1173, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100000100110011001101001011011001110110111111111000011111000010000100110110110100101111111111011011010001111001101000111010; 
out1174 = 128'b11100111001011100010001001100010011110011011111011010011001010010000010110100111110000110011000100001011010001111001111101010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1174[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1174, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011011110011110001111100101001011111011000111011111001111110000010101001110100100110001101000110000110010011100011000111010; 
out1175 = 128'b01011110011010110011011100010000100101000011110000011101100111010000000100000100000101001110010011011110011000000010111011010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1175[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1175, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100100111111110010000110011111011101100110001011000100011111111100110110110101001101001001100011000101011100001101011000101; 
out1176 = 128'b01101100110101111110000100100101110010010011011011100010110010110010101011100001000001010100111100110111111001011001010010010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1176[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1176, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100100111011011111011001110010100101010100010100011100101001100001010011101111111001000000011111111011101001110101110100000; 
out1177 = 128'b11010110011100001100101001000010111100000000110100111000101000000111101001110011000110111110010101010111000000111110100000010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1177[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1177, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011100010010011100001011001100100000011000010000111001101010001000101101111110011010000111111000100011100111111101001000000; 
out1178 = 128'b01001110010111001110001101000111011001111111111100000101101000111101011101001001110101101101010100001101110111110001000111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1178[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1178, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111010001100011000010101110010110000011000000011000001001010101010000111110010111110001010111010011100110000000110100110010; 
out1179 = 128'b10111101010011011101001011011101110000110001110011100110111101110100110110001100110110010111100111010101011011001001010110111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1179[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1179, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111011001010011100000100001110000111010101110000111001001010110101111010011011010100110101011010101010100011000110100011011; 
out1180 = 128'b00111111010010110011011000111000001100001010110001001011111011100011001100010011010100101101000011000010000110111001001110110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1180[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1180, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000110011001000000101000101011110001111101000011001100101100100011011110011000101101111000011001111011100110001110101100100; 
out1181 = 128'b01100001010000000110110001100011011111001000110111101000110110101001111100000110010100000100011111011111001000011010001011000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1181[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1181, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001000111001100001000100000011111101011111110001110010010110111000000011101000011101110011110101111100101110000000010011101010; 
out1182 = 128'b00010101100111001111001110110010111010010110100110000101010100000101100111101001101110111101111111101000010110101000110001110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1182[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1182, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110000010011111111111001011111001010010001010001101111001101100010101101111010101010010010111010110101010010110110100001110110; 
out1183 = 128'b01010100111000110001011101001000001100100011111000010011010011110110111111001010101111111011111000000011111110011001100001001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1183[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1183, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001100010000100101101110011100101011111100111001000100010000101010010101000110110001001100000111011001010100001010010010101; 
out1184 = 128'b10001001100110111000111110111111010101010001011001011101100010110000111001010010100010100000111001001011001101011000010111001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1184[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1184, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101101101010011001100001100001110111110110001101100011011100101000111011100000101110110110100001000000111000011000100000001; 
out1185 = 128'b10010001010000010000010001001000110000100011000011111000010011011111110011010010110100111010000000111111011010101000100100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1185[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1185, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000111111110110010110101110101011000100000101010111010110111110000001010100110110001100100010110101010011000111011111000000; 
out1186 = 128'b00000011000100001111010000000011010111010100101100100100011000000100011011110011000100001111010100000011111010010100110001110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1186[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1186, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011011011000110111110100100000110101000001111111010010101011011010111101100001011010011101111011111101111101100101100010011; 
out1187 = 128'b01000101000111110101011010010011000010001100010101100001001111110010010001111001111001011010000100111100100001011101000100100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1187[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1187, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000111010000000110101010101111100101111111100100000101110110110011010110000000100100011011011011111100001111010111001111001; 
out1188 = 128'b10000010011000110001100110011011001010001000001010011110000101000100101010011010101110110111000111001010110100010101000100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1188[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1188, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011111011100110001101101100110101010101011110110110010111001111011110100100010000001011100010000111010011111000110101000001101; 
out1189 = 128'b01100111100000010110101000001110100111010111101111100100001111110100111101111111111000110101001000001010100100110101010110101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1189[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1189, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000111010000100110110001101000000011010011011000101001101010100001011110001110011011011110110111000101000000000101001110111101; 
out1190 = 128'b11101101111010000110000101010100110011000010110000000110111011001011001100001001110111001010011001010110110001110110001000110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1190[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1190, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010001010100001000101110010010110100010100111100011001100101000110100001000000001001000010100110011101010110000101011100101; 
out1191 = 128'b00100100100110110100001101101011100111010100001011010111001010100101000100110110101010111101010111110010000010000111101101000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1191[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1191, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000110101001101111011110011001010010010010101000001001001100111011010101011010100010011001110101011110111011001000100111101; 
out1192 = 128'b00001000010001101011100101111110101101110001010110110110100010000000111110001111000001110001111111000011100101011110001010000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1192[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1192, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001011001001001100011111111110011111100000010110101011010110001101011001101000100001100001000101010001011101101110010001000; 
out1193 = 128'b11010001011101011011101110010000010101011000100000011100101011000101110100010011011000110000100000010010011001000010011101100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1193[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1193, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110000111011011010101010100100111000011001001110011010010110100010011100010111010001010011000110000101011001100101001101010; 
out1194 = 128'b11001111011110001101111011111000100001101010110000001010100010100110110010010111110010111100000110111110010011001111000100010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1194[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1194, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011101111111001100010001000100000000000100110010101010110001110101110011110011110100001001110110010000101001011111000100011; 
out1195 = 128'b00110010100101010100110101101110001110111101001001011001010000001100000100010111001100101100001011000101100101011011001001010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1195[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1195, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100111011100111010111100010101111010010100010000011000100111110011100110001111101000100111101110101011101010010011110011001; 
out1196 = 128'b00010110010000111110011110010100111111111110010000110111011100100101010100100001010001001101001111111111000001010011000001001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1196[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1196, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000011011111110001000011100111010111000000010101011111010110100110001111100100011011111110111101100010011011101100110001100; 
out1197 = 128'b01100101101010100101111101001100010010011110011001011110001010000100110111011010101001001110010001101111011110111111110101011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1197[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1197, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100101111111100111100001000011011111100010010011101101111001111010010011000010010000000000001111110000101101000100111100110001; 
out1198 = 128'b00001001111011100001101001000110101000111100111010110000010111110101011001011011000100111011011011100101101000010100100100110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1198[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1198, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010010000101110010011111101011001001101011111100000000101100101101100101001110010101111110110010111101000110111101111101011011; 
out1199 = 128'b10010010101000001100001010111010011111110001101010000100110000001111010110010100010110011101010100011001100011100111101100110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1199[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1199, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000010110000110000000001110100111000000000110100011100101010111001101011100000011111000000001000110101010011010110110011110; 
out1200 = 128'b11001010011110110001100110011010101011001111000100110100011110101100001011000010110011001011111111110100100011010100000000001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1200[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1200, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011101100001010101000101010000111001111101011100110000110010011000011100011000000101000010001010010110011011100111110101100; 
out1201 = 128'b11110110010110110111011111101011010000000011100001010111111110110110000100100110101010110001110111111111011001011010001100100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1201[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1201, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100001010111100010001011000110011111110001101100011100101001010000101000000110010100100001001010011010000110110100000111111; 
out1202 = 128'b11000000010011110101100101000001001010100011011001000111001011000010011101111101111101010101010001001010110010011011101011100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1202[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1202, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011001000001010001001000100010110101011101100010110011000001110111001001010111101100001110110000000000111010101111100110101; 
out1203 = 128'b01000111010110000110110100010010111110001011111100101110011010010001110011010001001111110010000001101001101001011101011011101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1203[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1203, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011000111100011101000111110110111011110000000011010001110001111101001000010111001010001100100101000101110001010111000011111; 
out1204 = 128'b00101111101101011000100100101001010011111110100001101101001100000110101110100010111011000110001110000100110000110110111100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1204[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1204, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101100010000000111100111100001101100001011101100100100011111001011111110101110010011111001010010100101111111000101001011001; 
out1205 = 128'b00010110011000101101100011111111010110000101001011001000010110010101001100001110001001111000101001011101010111111101010100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1205[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1205, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101001110000100010101000100111011011000111000000010100100100101100011110110111011111110001100100111000010101110100000001001; 
out1206 = 128'b00100100101010101101110111101001100011111011010100010011001010000111000110110101110010001110001011000110011011111100111100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1206[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1206, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101011111101000001000001010000000010100101001001011100011010110101110111110000111110111111011010010001111000110001101110100; 
out1207 = 128'b11111010000100111110001100111101101000110110010001100101001101100100101100001001010000001111010010110001010010110010110100001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1207[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1207, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010000000010010001000100101010001000010001111111011000000100110011100111010100111100000110101010001010110011010100000011000; 
out1208 = 128'b00110000001011010001000110110100110010111100011111110100000110001111000110000010010100000010001101011110110010101111100001110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1208[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1208, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001110010100101101110010000110001001011000001000000001101011010001011000110010111101000111100110010101000100110101011000001; 
out1209 = 128'b00011000000011100111101101111111001001001000010100010011101101001011110000011000010110011000100011010010101111101010010010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1209[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1209, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010011001011100101100011101101010110110010001000000001010001101000000000101001011010000011011011110101101010000011110111001100; 
out1210 = 128'b10110101010101011000011101111011100000101011011011000010010100010111111011010111101100101111000110000110011010100101000110110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1210[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1210, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100001000000110011011110111100100000000110000100111100010111010001001010000100111011101100001110000100000100110000010101000111; 
out1211 = 128'b11010000010110001001110001101000100000001101100100001100010000011110111000100101001011010100100111110111000011100110101011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1211[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1211, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010000001010010010110101110111110111110000110010100010011101110010001010011000000111111100011011001001110000000101101111110; 
out1212 = 128'b00111000011010101100110000110001110000000101011010001011000110011110000001101101111011110110110010010011101010101101011001000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1212[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1212, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011010010011110000001000000101011111100010001110010101000011001001110011101100011111010000110100010110001001010100000111001; 
out1213 = 128'b01101110000011111010111111101011010110101010101100111100001101111110000010111111111101011000101000001111100011110111100010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1213[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1213, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000111111010100100000001100011001010101111100100001100110111001001101110011110011010101101001001010001111011110110011100111; 
out1214 = 128'b00001110001111000011111111100001101111101101101001001001011110011011010011100110101000111100110110001001101000011010100000111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1214[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1214, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001101001010101111011110101011000111111100000110000110001000011101100011010110010001111011001001001110110010101101010100000; 
out1215 = 128'b00011000011011010100101111000110101001111010010100001011010000110100101011110011011110100010010011110100110111110001100010100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1215[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1215, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100001111010110001011101100110101000001001010001011000110110000010010010010101010010101011001110010011000101111101111110001; 
out1216 = 128'b00111010001000011110010110000010111100100100001000011011001100000000110010000100100110100110010001111011100001110001000110011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1216[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1216, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111100001110101011101101011010001111100110101100110001000111111000001101111000110010001011011101010100011000011101111011000; 
out1217 = 128'b01000101111010010110000100001001000001101111011001100110111000011001000010111010111111011001011001000001101000011111101110100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1217[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1217, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011010100110111001100001010011000100101100101001100100111011100101110000001000001000111000010110101000010001001111100010101001; 
out1218 = 128'b10000110111111110001111001100001010111100110100111001000000101110001011010010110001010111101011101110100101101001100110001011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1218[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1218, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101010111010010100101011001010010110100000010101010110011001100001010110000001110101010100000101100110001000101010100010101; 
out1219 = 128'b11100100010101001100110000001010100000110111111110101111010010100110011101101001101010000001100110110000101000111011001011101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1219[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1219, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011101100100100010001001011010100000000111111011101011111100010101100111011110110011010010001111000111010100011010101111011; 
out1220 = 128'b01111000100101101001010000010110010000111011101000000110101101110011100001101000111101010001011101110101010011011010111001111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1220[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1220, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110010010101011100110011110011100111111010011010010101100111001111001111011001100101100111001011011000010011100110001001110; 
out1221 = 128'b11011101111001110001001100111001100101001011110100001010101010001101011001111010000011001100011101011111010001011101110111011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1221[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1221, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000111101101000110100000100100000110011011110011001110111111101011000010100001001111010001100110001111001110111110111000010110; 
out1222 = 128'b10011011111010010011101011011100011110001101100110011001011101010000011101101111111101111100010011101111000001111000111110100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1222[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1222, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111100101100100011111101100011000001011111110001110101001001101001000001011011110001110010101111100100101010111101101100000; 
out1223 = 128'b10001010000110110001010111001000100101101101000101101100011100110111100011100111101100001111001011101000000010111001101000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1223[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1223, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110111001111000111110010100111000111010000111000111101111001100000011010000000101110100000110010101000001111111100101110100; 
out1224 = 128'b01110111111001101000101100101011010111000110111100101001111001110111101011111100001111011010011000110010110111011011101100010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1224[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1224, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111111101001000000101101101100100111111001110000000100000001111100011111011110000000111101111010101010011110001000111110001; 
out1225 = 128'b11010001101001100000001011010101011110110110011000101001010111111000101101010101000001010001010110110111011101111000111000110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1225[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1225, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111000011000001111100000110001010000000110000111000101101001001101000101100000101100000001110000000100100101011100001100100; 
out1226 = 128'b10000101011101010110100011001100001111001011000111010101101010100111010010010011101000011010001101101110001000010010011011001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1226[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1226, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001111111011111110001101010100100001000111011000110101000100101001100000010000111011111100011001111010101001101101010111010; 
out1227 = 128'b10110101010110000101010011111011000000000101111101011011101101001110110010110000110011011101010110010001000111111000011110111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1227[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1227, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001111110111100000001100011100110110110101011011001000010001010011100100101000011010111101011011100111010100011100001111001001; 
out1228 = 128'b10100001001101101011000011001010000101000011010010010001101110000111110110111010111100111110110111101111000001001011001000110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1228[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1228, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011100100100110111110000100100110000000110010110110000000101011100011110010101111110011110000001110111101100001001110000001; 
out1229 = 128'b01110011110000011011101010111111001000000111101110100000000111110010010010110001001100001101111101011111010000111100100011011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1229[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1229, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010001001101110110111111100000011000101000100111011111011111111001010100111001111100000110100011100010110000000011101111010; 
out1230 = 128'b10110010110111000100110010001110010101110011100000000110011110010110110111101000011001110111100010111110100010001101110011110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1230[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1230, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101100011111110111101010001001100010110000000110000000000100011000101100001110111100100100000101010000000010000010000110010; 
out1231 = 128'b11101011010101000000011001010000000101000011100100101110000101001010010101100011100011010011101011011000111000100000100100100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1231[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1231, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110011011101110111000101101011101001101111111101101000011100100101000010000000000011101001110100110001101001100111001001001011; 
out1232 = 128'b10001000111111000001011110110010000101110000111111010110010000010011100110010011000110011110100111000000000111010010001101010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1232[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1232, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000000100001001000100011011110010010011110000001111001010111010100111111011111100000011110101010000001010101101111111010111; 
out1233 = 128'b01110010101000010011100010111001010011001101001110010010110010000010111000001010111001111100111001001111110000111101010110111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1233[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1233, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100011010100101010011110010010010110101110001001111110011000100111010000010100001011000111011110100010000000100111011011111; 
out1234 = 128'b10011001111010101000010111110110011011000101110110010110111101000011011101000110101000011001111101111000110110011110110011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1234[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1234, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110010101011101101100100100000010011011010000000000011111000010101000011010001010001001101101000101010111111100000100001000; 
out1235 = 128'b00100100011110000001100000011101101110011100010001100000110001000000010101110000001111010011000001100010111101111110111011111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1235[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1235, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101011011001000101011000010111001010100000001010100110110010100010010110111100111000101010010111001100101111000100101000100; 
out1236 = 128'b10011000110010001000000100100000011011111111111010010110100101110010111101111110111100000010110100111000000011101110101000110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1236[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1236, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100011000000110110011111101101010010000001000000010110011100000111011000001101001001101111001101111111000001110001010011101; 
out1237 = 128'b11110011100000001001011110000011111111000011100001010010101001001101100110101110111100111110010101000011111001110011011100011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1237[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1237, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100001111110001111111001100001000100100000010011111110100111111100010100111001100110100001111110010100101010001010101011101; 
out1238 = 128'b00001001110000000001100110000000010101111100111011011001000101101000011100110000100111000010001001010001011100111101000100010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1238[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1238, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011001010011010010111101001001101001111010010001011011001101111001100101010001100111011010011100011000001111011000100011111; 
out1239 = 128'b01000010001101011110111101010000000100101111111100100110101011110111100001001001100110011111000011110101101110010101010100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1239[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1239, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110101011001000011110010000010001101001110010110000000110000011100011000011110010011011110110101010010111111011100101111110; 
out1240 = 128'b01101010110111000010101010000101001000100111111111000111010011000111001110101010111101010101001000111110011010111001011011000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1240[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1240, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001010101001101100100000010010011001101100011011110000010011010101000100011000110100110100110001001100001111011010010010000; 
out1241 = 128'b11111011100101100101100111010001100001111100111010001101000001100010000101001101100011001111111010010011011111110100101010000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1241[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1241, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101011101110100011100101110100101001100111001000000011111011101011111100000111001010000010100100110011110101001000111100110; 
out1242 = 128'b10111011100011110010111011111111110001010111111100111111001001110001110101101000000101010010111101100001000101100001000000001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1242[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1242, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001001001101000011011011001111011000100011100011011010101111011110010110101011000011100010011100111100110001110110001000000001; 
out1243 = 128'b11011000011000110001100011000110101011101100101001010010100101111100011010010000011001010001000000010001111000100110100111011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1243[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1243, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010000000010001110110000010110111110111111101011111001010010010110001101010101000110011001101001101100010010100101110101010; 
out1244 = 128'b01011111110010010000000001110011011000011111100110011001000111111001110011100010101110010010011101001011001110111101010111101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1244[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1244, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100100000111011010001100111010011100001101100001011000111010010001000010001010010101010010011110001101011010100010010010101; 
out1245 = 128'b11010111110110100101011110100110011101100100011001011010111010001001000110000000100010000100100101111111110111100001001110010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1245[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1245, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110111001000110000011110111000100101110111001010001001110101011000001101001010011001000100000100001100010100001001110100100; 
out1246 = 128'b10001011000100010110000000010011110110001010000011001001010000011011111100000101110010011110010001001001100001101100100101101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1246[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1246, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000000110001101010011100011000101100011111100100101010101100101001001110011101010110101011000001110101001011110011100111101; 
out1247 = 128'b00110010100101001100100011111100100000111010100000111100100101110000111000000111010001001110011110001001101101010011000000001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1247[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1247, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110101101111110110011101100011111011000011111000101000101111010001110111010001100010000000001001110110011000011010111010011; 
out1248 = 128'b00111110000010111101000111001010100110101111011001011101100101100100000110010101101111100100101000001001100101101100111011011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1248[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1248, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000110111000001000101111000111101110000111100111110111001101111001101101011001001110010001101000011101111001100010000101100; 
out1249 = 128'b00000011010111101000111100111001010010100110101110100001110111011100011010001001101110011010000001100001110100011111000100001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1249[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1249, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000001101010100111000000111110000110100101011101010000110001010001100011111111111011100010111011000001100111100001100101100; 
out1250 = 128'b10110110111010001010100111110000001001001100101000110111010100000110110111010110111110110100110000001101111011110111000011000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1250[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1250, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010000100101101001010001000010110000111010001101101110001011010010101011111110000111011101011010011001010010100100111011101; 
out1251 = 128'b10101000101101011011110011010110010000101110011010110001000101100100110001100110010000110111111111010100011100010000011000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1251[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1251, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010011011101101000100000000000011010011000000010010000011001100100100011101010010010001000111100000110100001100001100001110; 
out1252 = 128'b01111011111110000010011010100101100110101011111101001100110110100110111110111100110011101000110001001101101000101100111100110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1252[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1252, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011010101111010101000100000010010101111010000110111101100001101000100110100001001111111000100011100101001010010001110010101; 
out1253 = 128'b10111101111010100100000001100011110111011100011010100100010110111110000000001010001001100101001011101000100000010001000111100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1253[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1253, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101010001001010110100011110110101011100001110101001001011110111000000101100001010101010000111101110111100011010011001000011000; 
out1254 = 128'b00000011100111110110000011111001001100110001101101001000101000000001100111001011111101110000100100100000000010100011011011110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1254[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1254, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011101011100100100101010010001001111111001100100111011010001010101101010110010101110101110101111111101100000010110110110111; 
out1255 = 128'b00010010110000100101011000101111011110101110110001101111101101001000011100101111001010000101100011001100001101001000111111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1255[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1255, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110101000000110000100010101111111111010000110010101111111011010111100110010100100100100011000000110001010100000101010101000; 
out1256 = 128'b10001100000110011001010011110001110001111100000100000010011000100110001100001100010110011010010101000111100010100001000010100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1256[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1256, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111110110111000010111001010010111110000101101010000001110111010000100001101101110001011010000011001111010010010101010000010; 
out1257 = 128'b10101010110000110000110101100001111010001101100000001001010000101011010110000101000010011000111101110000110000111010101101010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1257[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1257, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011001000010000111111101101010001011000100001111010111000000101010100000101111010010010010000011000100010111111000011100000; 
out1258 = 128'b00011011001111100111101000101101011011100111101000011010110000110111101011000010111000010010011110111001001001100000100000011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1258[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1258, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010011001101010001001110111011000010111000110010001010100010101100010111000110001000111101000101100001010110101110110010011; 
out1259 = 128'b10110110100000011100101010010110110011011100111111100010001011011011111100001101111000101010110010110001101000111000011001001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1259[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1259, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110000111100001000100001101010110110001101111111011110001000111100100100010100001001101101101001011011011110011011011101011; 
out1260 = 128'b10001110101010010111101111110100011100000101111000100101111111000000100001100101100101011111000010100001010100010110000110110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1260[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1260, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000010011101101101110111100111011010001000000100000101000110111110101010101111110000111111101111010100010011100010001001111; 
out1261 = 128'b11001110111001000011111000011010000000100011010011000100010100000110110010111010100111110110111000101010100001011110010100110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1261[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1261, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111101110000111001110010111001111000111000001100010000000110000100110000010011101001111101011001101001111011101101000001110; 
out1262 = 128'b11001010010111011111001110010001110110001100100001011000101110101010000110100110001111111100110001110100011110010101110111011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1262[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1262, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011100111011110101101101010011110101101011011110011111001111010010110111111110000111101100110010010101101111100110100000110; 
out1263 = 128'b11011000100000010000001000000100010100111111001011010101010011111101010000101110101010101001110000011010000011011010001011111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1263[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1263, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000101111111111000101100000010110100001010011110011010001100010101111101010011111111001011101111011011011111010000110111011; 
out1264 = 128'b11111110101011011110101001010100101101100011000011000111101001011110011011010110111000111010000110101101010000001001100000111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1264[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1264, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010011110111000010010000110110100110001011100011110001100101000101000110001100001000000110001110101111001101110000010110001; 
out1265 = 128'b01110111111000111101111101100101010011100000001100110000111001010111000100110010100110110010110010010110010011100101000000101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1265[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1265, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011111110000000010100111111111011100011100011110111101110001110110110000110101000011111011110101000000101011000100001000101000; 
out1266 = 128'b10100101100011000101111011010011110010001010100111111011110011101101010010011010000110101011101100111101000110011101100010110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1266[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1266, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111110100000011111111101110000100011100000110110010001010101100000001001000000111010100000101001000110010000110010110010110; 
out1267 = 128'b01110001100100011100111111111111011110000101101100110011110001010101001101101111101101000110111001100100010110101010100000100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1267[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1267, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101100110001001000100010010010110101100110001010010001000110110000000110011111100101001001000001000100011011011111000110110; 
out1268 = 128'b10000101011000111101001111100000010100000010100011100000100111010100100011100100010010101101111111101110100100011000000011101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1268[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1268, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010011100011011100001000111000100010010100100011100010111010100010101110000110011010110010011000010000110011100011001110011; 
out1269 = 128'b11000011100001011100110111000001110000000001100100111010011101101100001101100000001100111110111010111101001100111110100001000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1269[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1269, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110100111110110010101110101000010101100000101010100110010100000001110100010111101111011100101111001111011010100101100010010; 
out1270 = 128'b10100100010111010111110010000100110111010100000101000001101100011110000010111010110100110000100111011100100010101110010000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1270[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1270, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011100000011011001001101110110101001000011101011010011100011001011100001001010000000111110100100000010010011000011010011110; 
out1271 = 128'b00111011000100110100111110000100111010000111111011101111010001110001110010010001101101001010100100101111111010000111111000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1271[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1271, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011010100111111001111100101011001110100001100001100101101110011101010010110010000001110011010100001010110101010011110010101010; 
out1272 = 128'b10010111001011011010010111000110010010111101101101110011110010111100011101000011010111001001101010111110101000101101001011110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1272[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1272, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010111000100110011010101001010111111010110000000000000110000010000001111001010011001010101100011011000101101111100001101111; 
out1273 = 128'b01100101101110100001011000010111110001001111111100010100000101111101100110000111010010010011011111010110110001001101010101110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1273[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1273, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111000111000111110101001001100011101110000001100010010010111110000110100011111000001001101111110101110100101111000000001111; 
out1274 = 128'b00100001010101001001010110011111011111000111111100001000001100100000000000000111100010111111011000110000100010101000000100010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1274[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1274, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010111100100000111111000100011111100110001001001110011010100100111111001001100111001100111111101010100010001100001011011010; 
out1275 = 128'b01011010010101011110000110001011001110110011001100101011100010111011100101000010111110100001010010011101100011000110100110110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1275[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1275, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001010111001101100000101001111100100010111010111000100011001011111001101010010000011010000101100001111001001001100101000100; 
out1276 = 128'b00010000111001010000100010101000010011111101010001000110000101010110011100110100000111100111001100100111011011001011010100000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1276[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1276, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101101011000111101110001110011000111010011001000110011101001111101110100011101000110100010110011111011111010101110100001000; 
out1277 = 128'b10110010000111111100100010011010001011010010100011110011110100001001001001111101000101101010111001010101111110101111010000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1277[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1277, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010010011110010010010011111101111110101100110011001101001000110111110001101110110110110101010110010001101111110100111100011; 
out1278 = 128'b00101011111101100100110010010011001111000110100101010110000000100011100111111000110010110100011000000110001001111100011101101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1278[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1278, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101001000110110111000111000010010000101100010010011011000010100110110000001100000110000100110010000111110010000100100101011; 
out1279 = 128'b10110101100001010010100010000000101011110000010100100000100011100011001110111000001110110001000100000010001000011110110000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1279[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1279, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000010001000001110101011111001001001101110010100001010010000000010001000111001000000100110001000010111101011010010101111100; 
out1280 = 128'b11110101000100111001010011001011011101010101010110100010001011001010011011010001001010100101010001010111011010010000001111100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1280[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1280, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011010111101011011001000110111100111011111010100010011110110110001100111010111001111101000010100111111101111000110100001100; 
out1281 = 128'b00101101101101001001011101111101001010000001010110010100101001110100111011101100101111011011010000000111010101110101001110100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1281[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1281, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001101110110011000001100010101111011111110100010011011011100001111101111101001001000001101101101011000101110000011100001000; 
out1282 = 128'b01011111000011101011111010001011000000001010001010011111111011100101101101000001001100000110101011011111100100101101110110111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1282[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1282, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100000101010000101101100101010000101101010000111101000011100101000010111100010101101001100000010010010100000000000011000111; 
out1283 = 128'b10001100110110101000111100001000011101100101111000110110011100000100111011001000001101000110000110101000011010010001100011100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1283[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1283, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001100010101001001001001010101110110101000001000110100010001101100100111111111001001101011010011011100000010000000100111011; 
out1284 = 128'b11111000110111110101100000011101111100101101110101111110010000001111000011011000010100011011100100001101001110000001111101000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1284[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1284, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001001011011100111010000001010101001000000100010011011111000000011100101010000010101101001100001001010001110000100011111010; 
out1285 = 128'b01010101101100101001100100101101101001011100010100001111100011101001110110000001101010101101100101100100010101101110000111111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1285[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1285, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011001110001001111101101100001101111001111011011100101001011100111001011000101101100110001011000100110111101000000000101110; 
out1286 = 128'b10110011101011001000100001000001110100101010110001101010000011111101110001011101011000100111010101011101010110011001100010111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1286[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1286, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010010101000101000011000010101001100101111111101110110011011100111000100110100100101010010100111101101011001101100101010001; 
out1287 = 128'b00010000101110111101101011100110101000000111100111101011011010111101100010011000001100111011101111101000111111001110100101010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1287[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1287, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100111110010110111100001011110001101000010011100110100100111100000111010101010110001111100101011011101000011111100110110000; 
out1288 = 128'b01000101001001100010111001010111011010111011011100011110100011000100011111001100000011000001010101111111101001001100010001001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1288[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1288, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111101111001101010011100101001010011010101101000111101001011111100001110111110100111111001101001011111010110110100100000010; 
out1289 = 128'b10111011000000001011010010010110110000111101011111001000011001111111010000001100101101010101100100000010010000000110111010110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1289[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1289, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011100001110110000011000000001011110001100101001100001100100011111010000110001011110110111110010110101000011100101011100100; 
out1290 = 128'b01110011110111110010010011010010111110001001001111010011111110010000001100010100001101001001001010100010101111011110010001111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1290[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1290, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000010101110101010101001100100100011011001100011111011100101001001001101100001011110100101101010101100001011110111111000011; 
out1291 = 128'b10100111000000010010010010110001111010011010111100010011001011101010110001101111101001110010110000001001010000101110010101110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1291[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1291, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000110000100011001011011101000011100001100011001111001011000011111110100010011110011000101110100011111101000100100100000011; 
out1292 = 128'b11111111001001101111110001100000011100001111001101110010010010110110011111110101000000101011101100001100111001000011001111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1292[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1292, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001101111011011010101010001011011100011001111001001010011101011101110110000010000010101101111110111111110011111110010111101; 
out1293 = 128'b01100001111111100110010111100011011110001110101101000000110001110101110100101111011011001100011100110110010001010001111011010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1293[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1293, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111110000111011000101001010011111100100110101100111101000010011100010001100111101001101001000011001110010010110000011010000101; 
out1294 = 128'b10101011001101001001101001001000101010101010101101111111110000101011001100101001101011101111001010110100100100001111011000111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1294[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1294, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001101011101101011001110011111010111100111011100110010001010101101011011110000000001101000101111001000001000110011001110100; 
out1295 = 128'b00011000000101001110110000100101110110101001011111011111000111110101010110011101101110101101110110111001101111000011110010011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1295[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1295, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001011010101111110000100100010001001101010001111101101110011111101001000010000110000001101001101001001000110111111001010001101; 
out1296 = 128'b00011011010110011000010101011111010001011111100011111100000010110110100111111000001000101100100101100010001000011011100011111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1296[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1296, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110011101001110010111101000000011010011001010001000000011000000101101100010001101100010100111011010101111111101010000010011; 
out1297 = 128'b01111001010001100100110011001000011001100000000000111000000111110100111001111010001111011101001111101110100001100101001011110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1297[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1297, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000110010010011000100110110110000010011001000010111011100000110000110011110000011000000010000110100100101110001101001001011; 
out1298 = 128'b01010101111011100000010011100110011111001001110110000010100111101101001101101110001100010000010110111010100011101011100101111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1298[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1298, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101101111111011101010101101101001100101101000000000000011001001101100100110000010111101101000000100000111010000000110010110010; 
out1299 = 128'b01100101110000110111010101001001010100111010111100100011111110000001111110110001100011110111001101011000000111000011110010100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1299[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1299, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100111111010011101011100111000011001110011110111111101111110111010000000000100001100001011101011000001101010001001111010001; 
out1300 = 128'b00101110110010001101111111010001001111110011100000000110001100110000001001100100100110100100010101111100011001111001100000000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1300[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1300, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000011000100001010101011001100100111101110001010111111001101111010110101101010101001010110110110011111000001100011110101001; 
out1301 = 128'b11100100100111111110001101011010111010000000100101110001110001011000110100001010100001101110000111011100100010000110101111101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1301[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1301, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101100100111011011010000101000110001001010000000010101101100011100000111001000101100010100001100011101100100000000111110000; 
out1302 = 128'b01000100000100011000000000010000001100011011001111110011110101000011010011011110000110001001101000111101010010110011101100110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1302[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1302, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010001111001001001011000110111000101000010101110101001111000010011001100010010101111111111001000101101001110010000111110101; 
out1303 = 128'b00010001000101011001001001101000111011001100111100001011011101011001100111111111110110101001011100000111000100100111011001110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1303[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1303, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010100110011000110010001111010010101110001011010001010011011000011000011001110111100100001101100001011111001111110101001000; 
out1304 = 128'b10000111100010000101000111011011110101010001110011001101111101101000111001101000000111000111000010010101111001110000111101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1304[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1304, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100001010101110000010100001011110010110000000100110010001011011001101100001011111000111111100100010011101001000111110110000; 
out1305 = 128'b10111011110101101000101011000100101001111111011101010111110101110000101010011001010010101100110100101100101011111111100010010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1305[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1305, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111101110101000110001101100010111000101000110000011111100100101100110000010011010101000001101110111101010011011110100001100; 
out1306 = 128'b00110001001000001010010111111100011110001011101001100110101111000100010111000101100110001100001010011010000001101000010010101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1306[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1306, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011000100001001111110011011111010100100000111010010000011111110011101110101100000011101011110011010010111010110000010000000; 
out1307 = 128'b10110101111111101001111001110110011111000111100101000011101101011001110101111000111000101101110110110001110000111000111010000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1307[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1307, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111001111010100001100110001011011101101111101000101110001110001110100000100100011110111101111000000100101000000111101000101; 
out1308 = 128'b10000100111011000100111000011111011110110101010100110111001001100101001000011100100101001111011011111101000010100101101011110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1308[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1308, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110110101010000101100100000010001100000011000100100101001011001010010101111101011101000101001101100010001010101101001001011; 
out1309 = 128'b10111111111000100000100101111110101001111000000001000101011000000101011111101101010100111110100010100011000101001100111100000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1309[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1309, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000110100010000110111001111100010011101011000101001110111000111111010100111010101111011110100011110000001000110000110110001; 
out1310 = 128'b11010011100100001011100101101101011000011011011010001101011101100010101011000110100010010111100010000001011000011101001101111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1310[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1310, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000011001110111001011011000111000000011110001101111111110000111101010010001011111001101111110011101100111110011111011101100; 
out1311 = 128'b10000101011100010011011110010000110100110100110011011010010111111101011010011000011110011111101100101010100101001100010101100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1311[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1311, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010000000110000100101001010110110001111100001111000100100111000000101100011001111011010111011110000010110000000111101001000; 
out1312 = 128'b10001110110011101111101100000110100100100110010110011000101101001001011011100011000000111010110110110001000100001000101010100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1312[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1312, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101101010010110101011001001000001000110001001111001110011001100110110011110111001010110111101010000001101100111011001100110; 
out1313 = 128'b01110100100001110101001101000111010110001101010100001111010011110010100111110011100001101110111010111101001111101010111101001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1313[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1313, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110101100111000001010101100111010000001110001110101010101100001010001011100100010001101101001010001010001010110110010110000; 
out1314 = 128'b00111001001110011111000101010001101110111010001101101011111100101001010001110110010011010110011111010000110000111100010010001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1314[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1314, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011100000100111010110101000110100110001100110000110111010111101110010101111011000011001101111110010010000000100001111111100; 
out1315 = 128'b01101000111110001111011010110011001111011101110100001111110001101110001000110010010111111000010010000101101010101100011111101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1315[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1315, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011110111101010101001001101101000000000000011110100100001001010000011001001011111101111011100001110010011011111000000011001; 
out1316 = 128'b01000101010100111111101101101100101010100011101111000100111101011001110110101100100011110101010100111011111101101111110101111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1316[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1316, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000010001001001100010011000000010010001110010111001111010010101001100110100011000101101111111110011101110111101100111101010001; 
out1317 = 128'b00100011111101111011000110000010000100101111001100111111000010111000101011000100100010101110011001110010110011010111110010101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1317[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1317, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100101111100100001000011000110010010010100000110010101000111110001000110011110001101110000010001111011000101101011111001101; 
out1318 = 128'b01010011000011110001001110111000011010111010011001010110001110011111001010111101010000001001110010010001011000000011110111000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1318[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1318, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111111110001100111100110101101110101111011000001110110110101011001010010000001111100101010011011011010001001001111101110010; 
out1319 = 128'b00100011001101000101101110011010111010000001101110010100100111001110010001111010001100011010110111111010100101101101100011101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1319[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1319, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011000000010001010100101101001011110110111100111111100010100011001011101011110101101011101111111100001110101101001100111011; 
out1320 = 128'b00101010100011100101111111000100000100000000100010110111010110011000000101111110101101010011111111011111000101001110100010001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1320[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1320, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001000010110000111001010111110000100011010011011010011110011011010001110100111101000111000010010110001101000001010011110011; 
out1321 = 128'b00111000111000100001010010011000000001110100010100000110001010100001010000111110101100010110100100011100011010000110101110011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1321[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1321, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111110110101000101001100011100110100111100100000001100111011010100110110001100011000101010100010101111100011011111100010000; 
out1322 = 128'b00001101010011101101000010011110111010000000101101111010110100000011100000101101100010100001110101111100111100001100111010011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1322[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1322, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111111110011000010011001100100100101000010011111101001101000011011111100110001111110001100110001111000100111010111101001100; 
out1323 = 128'b11100011111011111011101111110111110000000010001110110011111001100000001000101010011000110100110101010110101101100111101111110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1323[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1323, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011101001100111110000000010011101001010001011010011101000001101011110100001111101110101111101110010010011000001001000011001; 
out1324 = 128'b11010000111110100010000010001000000101011010011111100101101111111000011101001011011101111100010000001100100001011010111000011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1324[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1324, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010001100011011000000110101010111101011011010010100011001110010011111100110110110111100011011110011001110010001110100100000; 
out1325 = 128'b00001010111011000100111111110111100100000111000011101000010001101010010111111110110111000110110110101011001111110001011000000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1325[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1325, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101011010110000111111110110100111001001001101101100011110001110101101001001000100111010111101101000001010010111101110010101010; 
out1326 = 128'b01001110011111111111101101001000110100000111110000001101011010010000010001011000011000011111110011001101001100011001011001110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1326[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1326, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110100010001011100111100111100101110101010000100110010101000100011010000111111000011010011001111011110000011101111011111000; 
out1327 = 128'b11000100001001110100011001111100111001111110000100101100101001011010000001111011100011001111010101010001101111000111110101011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1327[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1327, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011101101111111011010100000011111111000000101110001111011010011110000011011111101011001110000100000101100111111100000100111110; 
out1328 = 128'b11000110110001001110010011010010011101000110010000001001100111111111100110110111000001110010101000010110100100110001110011110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1328[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1328, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111100000010011111011001010100000100001010110100010011000101110000001110101000000100101100110001100001011101111111110111100; 
out1329 = 128'b00000010001111111111011000111000010111110110010011011000101010101000010000111000110001100101011011001100110000111100111001101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1329[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1329, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011001110101101001010110011001101010110010100010100010010011000000110000010100110100111101101111010100100001000000100101101; 
out1330 = 128'b00100100101000101011101000011110111111100011000110011110111101000011010101100111100001000000111010000100010100101011010010010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1330[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1330, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011001100011010100000101000000010000000001110101011100000001100000111101101000100010100111111110011101001001101100000000110; 
out1331 = 128'b00100101100101001101000011100100000111000111101110111001101101000111000010001111100101001010111000110100000100101110101011000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1331[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1331, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100101111101000110001111011001010011010111010101001101011100010011110101101010011111111000011011001100010110001111100000111; 
out1332 = 128'b00001111011011011100100110110111100000000000100110011111000001111010100010010001001100111101110111001010110101111111100001001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1332[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1332, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110111110100011011000011111101110101001001101010011010010010000010100000000111000011010001101101100001110000011000110001110; 
out1333 = 128'b10101100011001000000100001001001101101010110110000111100010010010001100111111011110011110011111101110001010001111001110001110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1333[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1333, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110100001111111000011000011111001011001101000101110101000101011100010110010100011010010010010111100011101110111000111101110; 
out1334 = 128'b11001110111111010010110011000100110111100000100010010010010100100100111111111001010110001000101001101000111000011101010101101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1334[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1334, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000100001110000000011000000010100111011000101101111100011101010111001101100101010010000100111000101010011111001101001111001; 
out1335 = 128'b11101111110010101101001110010010001000001001100110100000111111111001010100100110001010011100111101011001110011000010111000101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1335[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1335, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111001000011010101111001110011001010100010110010110011110010110110100001010011011101011111111001101101001101100100111010011111; 
out1336 = 128'b00011110000101000110010011010110111001100010010010010111011111001000001010110010011001011100111001111110101100011000000110001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1336[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1336, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101111110010110010000011111101111011101111110010100101100111111001010111010001001111001000001110011101000011111110101101110; 
out1337 = 128'b00110100011100001000100101100101110011101110011011111000111011101011000010100010001010101000010100110111000101111010101101101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1337[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1337, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110000100011010011111110011111111010111111001111011001010110110000100001010001110111011001101001010001001000110010001011110; 
out1338 = 128'b01110100111100001010011110110111010011100101100110100001001111000101101011110110010011001000100101010011101110111101100101100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1338[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1338, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110111001101011100000001111100101011111110000111000010010011010010111110100000010011000010000100100101011100000011011101000; 
out1339 = 128'b10000101000111100100100100111111010101001001100111010001010111110111010001111001001000100000000010100001000010001011110001001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1339[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1339, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101110101101101010110100001110000101101100011111100100000001001111000011001011011101101000001011001111110110101011000000100; 
out1340 = 128'b01101111111010011000110001111000110001111110110100110111000001110000010011011110110100111100100110010101001000000110101000111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1340[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1340, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100111100101100111111001110111100000001100011101100101001001011111101101101000011100101010101001000011010000110110111000011; 
out1341 = 128'b00001001010100011110000010011001110100100100000101101001101101101110011110110100110111001101110011100001000011000111101100010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1341[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1341, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101001010000111111001011101010000101100111000000010101100011111100110000111110100000101011000001001101100100100000011101111; 
out1342 = 128'b00011101110010110100110001111110111000011011110010011000001100010110011000101100110000001010110010011101100000000101010111001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1342[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1342, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011111101111001110101001010000001001100110100011001010011111000001000101110100000011111110101001010111001110100011001110011; 
out1343 = 128'b01010100011001001001011111001110000100101101010100011100110000111000100010001111100101001001100010100101111011100110011110101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1343[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1343, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110010000101100101100000100101100000100000001010100111011000100111000111100011101111011101000110000111011101110010110101100; 
out1344 = 128'b01000000001110001011011111010100010000001100100110001100010010110110101111010011100000110011011110001001011011100011111101100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1344[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1344, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100110001100111000011000000011011101101000010010101111101011011011110111000011100000011011000111111010011001111101110100011; 
out1345 = 128'b11001101111010100000000101101110101100111010011000011100010000010101001011110110000010001001111100100100111101110111010010110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1345[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1345, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011000011000101111001011011111100001001001111000001110111111000100000101111110000010011011000010001000100111111010001010111; 
out1346 = 128'b10101000000100001110011111101100110111000110101010111111010010100011011110111101100101111111111100011101101110101100000100101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1346[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1346, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000111010001010001011011111000000000000101011010110011101010100001100011110011011111000011100001011100001110011011000101111; 
out1347 = 128'b11100110111011111101110000101111000001011100011101011001101100010101110101000000000101101101011100010001110001100100001010100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1347[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1347, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010000101101111111100100000011011110110101010101000010110111100111011111011110001000011010011000001100010110101110111001110; 
out1348 = 128'b01011101001000010001000001010011000001110011101000001010101011000001110110110101000011111101010101101000000111111111111100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1348[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1348, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011101011010100110100101011100010110010101011101011111000111010000100001000011110101010010000001001100111111101111110010000; 
out1349 = 128'b01101011011101100110001110101101100101110111010100110101001101101111110011111111101111010110110001000101101010110001000010011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1349[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1349, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010100100101111011010111000011001100100010111101011010111100111000110000100001011000011100101110101011001101000000000011001; 
out1350 = 128'b10010110001011000001011100101001000111110010100010100011110111101010111000110000111011011011000010001011110101111111110101001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1350[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1350, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101011110010011011101001101110000110101001010010001110111001101111100010000011111110011010110110001110000111010110100011111; 
out1351 = 128'b00011111001000100100000111110100011111101110100110101011111011010010011000111000101011101111111001101101000001111110100110010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1351[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1351, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101110011110001111100101101001011100000010001011111000001000010000111110111011001010000110110111010111011110111101000101001; 
out1352 = 128'b10100101111111111001011100001001011100001010100000100000100100110001110100110110001110000011101000001001101110010100001110110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1352[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1352, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000110100011100000001110110110110010111110110011011000101001010101100000101100111010111010111101001110111001010101000000000; 
out1353 = 128'b00010001011101000100101110001001110000011100111001100111010000110100100111001001101101101011010010011010001001100101110100000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1353[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1353, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001100101010010101010000011010100100011100110111010101010100100111111111001100111001111001100001011100111111010011010110101; 
out1354 = 128'b10101010001001101010001001101111011000111101000011111101001110000101111111001000001011000100010010100011100000110011101110111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1354[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1354, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000010011110100100000011011110010100000010000001111110001101000001010000010000100101000010011001001110000001111111011100110; 
out1355 = 128'b01010110111001001110010111001001011011100101101111001000111111011001100001110010111110000001001001111111101101011110111101010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1355[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1355, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110010100110011011000000111010100101100011010100010001010110111000101100111001001111000000001101101111110001001000000101110; 
out1356 = 128'b01011010011110000110110100010011101011100001010100000101110000111110011110110000000110010100001101100100010101011011000110101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1356[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1356, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010011110010110001111001111100101010101001101011000110011101101111001001101101011011111100010001010000010100000110101011100000; 
out1357 = 128'b00001001000010110101101110111010011101101101011000001100001011010100101100100111000111010110100001111110011101111111011011010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1357[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1357, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010100000001000111100010001110010001100100100010111110101111100001000111000000100110110010101111001110111000101000101000011; 
out1358 = 128'b00000100101110110001001111101101100011001011010110001010100100000111010010101011111111100001011101110100100111011011111011000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1358[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1358, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010000100111010110100101001100000110110000011001001110000010110100111110111111001110100001110010011101100010001001100110000; 
out1359 = 128'b01001010001100000111101111110000001010111001011111100011101001000110100010100100011111001000100101100100010111000101101011000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1359[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1359, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000111000010011111100010010010111110110101101101110010110110101010100001111111101101000001001101010110010100010100100001001111; 
out1360 = 128'b11010100111111001011010010000010101101010001001001010101110101111000111111110111000111001100000011110100001000010111001101010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1360[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1360, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100000101111011011000001101010111101010011101011011010110010000001010111100000110100001101001011001010001111100011100001000011; 
out1361 = 128'b10000100010101101100101111111111000110101100111000011010010001001100000110111100110111010100011010100011011110001001011010001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1361[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1361, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101010100011101011111101000010100111010100000010011000000011010001111010011110111111110101000110000011101010101001101111111010; 
out1362 = 128'b11100111111100001000000110100011000110010000100010000000101010110100111011110101010011101010000110001100111101000000110010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1362[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1362, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111001110000010110001111111100000011010000011111011001001010110111110010111101010001001110010010101111101111001111111001101; 
out1363 = 128'b11010001001101111001010011110000101101011000011101000110001101100001000100101000000100000111100001001101000000010000000110011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1363[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1363, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101010010000110100001001001000100101110011101001010111001000011011010100010000100001001111110100101100100100000100011111101011; 
out1364 = 128'b10101001011100110000111000000100110011100000001001001110101001111001000111111001010010101101101001011011011001000101111011110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1364[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1364, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011000101001010010111110000010011000000101101101011101101110111001010110000011110101100111111001000011100110010011000011111; 
out1365 = 128'b11011001110001101000101101000100101111100011101111010011100000000101000100010010101000111001011110000111110001011110000111111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1365[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1365, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101100111101100101111101001000110011100010101011000100100011011011100100001001010111011001110110110011011000111101111011110; 
out1366 = 128'b11001101000101110100100100100111110000011010011001111101000000100011010011010000010111000111001011101011011111011001110100000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1366[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1366, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111001111100010001010101111011011110010110010011101001000000001111100100010100101100000110111111100100110001100100011100001; 
out1367 = 128'b00101111111110010001011111110101111100111011001001011010101010111010110101110010100111111101010011110110011001110101000010000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1367[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1367, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000001111000100000001011000110010100000010010111101001001100111111110111001001001001011101010000001000000011000100101000101; 
out1368 = 128'b00110000101100000110110011110001110000010001011110110100011111011011000001101011001001000100100110011100001100011100001001111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1368[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1368, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000000111000000111000100001010000100011010101001010110110010100110001010010111111001111111010010011111110001111110110001111; 
out1369 = 128'b00000000010001110110100111011011001010010001111011100110110111011010000000010111110110111010010010001000110111111101101000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1369[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1369, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110000101100111011000010100100110110101010000100001111110110110001000000011011100110011000010011100110111110100100101110000; 
out1370 = 128'b01011001011111010100100100011100100101010011111000011000011000010011110101111110011111000010110110011111111111111011100010010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1370[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1370, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011101011110000110110010110010001010110101000011101011011010010110011101000000000110100011011100110110011110101001010111001110; 
out1371 = 128'b10000101010101111101101010010101111011011101101111001111111101101000010001101101011110100011110011010010111110000101010101110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1371[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1371, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010101000001100101101001101010001101011111011100010111101101010011101110100001000011000010100111110110101001101000001001111; 
out1372 = 128'b10000101010111010000100110100001100001110101010011111001110101001101111001110111101010110101001000001101110101100010110010001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1372[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1372, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100011100100111100010001011111001001110111001011101100000101000101110100101101101110000000000011101010010101111110110101001110; 
out1373 = 128'b01111111000100010000000110111111011101011100000000100010011011101001111010111011001011010010110100011101101111011011110100011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1373[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1373, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111001010001111111011001110101010010111010100101111100010100000000101001001110010010111010101001100000100110010111111110001; 
out1374 = 128'b01111111101101000111111100100010100100101011101010111011000000011110000101000000100011101011101011100110101101111000001011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1374[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1374, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101111100100010100100101000111111000110011101111001100101101010001100000101001010111010111010011010011111110001100100111001; 
out1375 = 128'b00001000101111101000011100010100111101011110100100001100010110110010011000110010011011001000010100110011001000101101101010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1375[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1375, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000111110000101000101100110110100100110110000011001111101001000111100101100100000011100001100010000000011000111010110111111; 
out1376 = 128'b01001001011010000000101111010000111110110110101111000010110110001111101001011100100111100100110110111010000001011101111110100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1376[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1376, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101110100010100111110101101110101110101001100000000001011000011111011110100100101010000010001000101101001001000111011111100; 
out1377 = 128'b10111111011110001101111010111000010101011100011111100011010000110000101100001110011111100111101101111110110110011010000011010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1377[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1377, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011000001011100110100010011010001101001001000010011011010100111100111101000101111011001101011010011100100100110011101000101; 
out1378 = 128'b10111110001100100001000110111011001111100110001010011111110101100001111110110001010110010110010110000001011000100101001101100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1378[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1378, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011010010110100111101000100110111100110101111010110111011000110000100111101010101100010000011110001011011111010111010010001; 
out1379 = 128'b11001110100111100001001101101101011111101110111100111111101010100010111111011111000001101010010011110010001100011000100110100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1379[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1379, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000100101101010110011000000000110111011100001000100000100110011110101110011100111001001101101001001101011110101010011000010; 
out1380 = 128'b11110011110110011111111101000110111001111110000011011111010010000111010000000011110000100001111001001110001011111001011001011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1380[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1380, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001101001001000000101000011010000110110111100011001010100100001101011101000000111011001101100110010100000100010101001011010101; 
out1381 = 128'b01000101000000101111110111000111101101100110001001000001111100011110010101001011011001001101011101011000011100100000010110100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1381[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1381, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110111100001101101110100001011101001011000110000001100011111010011111001101101000000110100001110000010011100000110010111000; 
out1382 = 128'b11010111011010010101001101011100001001110101111000001100100010100101100111100011010011101111010111001100000000110111111111101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1382[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1382, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010011101110101111000111111100101000000110100100000011000111001100000000100111010100011000001101101110101110010101111000101; 
out1383 = 128'b01000010101010010101110000110110000010010111110000110001001111001101001110010101100110101110110110101001111111011011011110001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1383[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1383, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100110001010010010001111110000011100100011011010011110110010000111000000000111110100001111111001111100111010001101010001110; 
out1384 = 128'b11011101011101110100010110011101110000101101000011001110001001010011111110010010101010100100011000100100000101011100111101000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1384[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1384, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110100010110001010111100000100000010010011110111100110111011110011001010110011000110101101101100001101111100101001001010100; 
out1385 = 128'b10010000001111001100101100001101111110101110010011010000000101010001100100001000110011000010000100110100110001111001110111101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1385[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1385, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001001000000110001011111001001110000011011110000000010110011000010111000111110110000010101011001100111110110001110100110000; 
out1386 = 128'b11010101100000101010111011101101011100010111010101011111001011011011000101011111001110111010101001101110010110001100010111111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1386[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1386, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001110010100101010101001110110000000011001001010110111010001111011111001110011101011100110001101001111011011010110000110111; 
out1387 = 128'b00101000101010000011000110101001110010001101011001101100101101111001010000100010010011111011001011001110011111011011110001110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1387[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1387, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010110101000100100110000100100010101010001100101011110000011100010010000110001000110010011110000011010010100111111001010101111; 
out1388 = 128'b10110100111011100101101011101110111100010101001110101001001011110001101111010010000101011011111111000000001111101111100011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1388[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1388, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001011011001010100000111001001111000101000001001100100100110001100011011011100100100011001000111111001101000001011010010110; 
out1389 = 128'b01010110001000101110011110010000010111011000111101101001110011101011110011101011110000010000100010101001010000010000100010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1389[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1389, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100000111010111001100001101001011010010001000011001001011011101100100010100000100000000011001010011100110011010101011101110; 
out1390 = 128'b10000010100101101011101100011001010101101100111110110100111010110011100110100010111001111100010001110010100000000100011110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1390[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1390, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010011010010111000100000111001001110000010000010011011100110100100000000100110000101110000000011010101011001100111110011000; 
out1391 = 128'b00011010100000001010111111011111110011100000111001010101011101001110101111110001111000000001110111101111011001101001010100010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1391[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1391, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111101100011000010100011100001101100001100000111011011101101111110001111010101001011111001001101101100010010010110110101110; 
out1392 = 128'b00111110001101010101100110011011101010111110000001101100101110101101011001111111011001001000010100100001001100100101100000000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1392[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1392, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001010101011101000001110001011011101110011010010101010110010110100001001011111100000111101110011001000101010010111100001100; 
out1393 = 128'b01110001000100011000010011110110010111010000100101000000000011100101101101011011101001001110001110011010101100010110011000110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1393[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1393, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100110001100111101001010011010111110100111101111101001001000110100111101001001001111000100100111101011100001101000010000111; 
out1394 = 128'b10000100000001111111111101010100110011000110110011101000100000101001001011110111111101110100111100010100011101111001001001110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1394[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1394, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010100000101111010001111000101111000101110101001010111011001101101010001001101010001100001001100000110011110110000010011101; 
out1395 = 128'b10101010010110100110001010000101011101111110000001100000000111011111011010100100100100011011100010000111100101110000101000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1395[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1395, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110001101111001100001011001101001100010011110110000111011111100001010010111101100001011101011011001111110011110101011000100; 
out1396 = 128'b11100011101011000010111110011010000101111000111100110100010001111010110000000101100100111101000000000000100101000100110001101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1396[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1396, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000100101001001000001100000100000100011010000111010011000111000100001101011011001010110110010110011110110000001000100101101; 
out1397 = 128'b01100101001110001000100100000111101011010010111101001111011001100110100111101101000000101101011101100110000101010111010000011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1397[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1397, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000100010110001011000000110001000011100010011011010101100011011100010010011100000010011101010101011001111100001000011101000; 
out1398 = 128'b11011000000100111100001100101001111100100010000011000010101000110101110100111110000000101011011101101111101110000101111100111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1398[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1398, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101101100101011000001100001101000011011010111100101000001001110100101101000001111000000101101001010010111011011100001010000; 
out1399 = 128'b01100110101001101100111101111011101111001100010001110111110000100111111010100001011110011010000101100110011000111011010100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1399[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1399, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111111001001100100000110111010111100010001101001000000001001110110000111110101110000001111110010111000111100000101110110100; 
out1400 = 128'b00001010110111001000111001001001111000010010000110001000011111001100001110000011011011111011010010101010001111101111010111010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1400[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1400, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010010111000010110010011011001101001001110001010110010101100111100111100001110011110010111110111110111011111010111011111111110; 
out1401 = 128'b01101110100100011001011101000110101111110000111100001010010100000111000111001101001100001111110000001101101110111001001111101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1401[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1401, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001101101010110010110000100101101000001111110010110110011000011101001111100110110001011100010100010011001011111010011111010; 
out1402 = 128'b11101110101011000011101110111111000101101100101101010110100111110011100110110111101000100101000100000101101010000011100100011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1402[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1402, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000111011000000011010000010111001000011110111100010001100101010101001010110110001010010011010111000110011000101000100101111; 
out1403 = 128'b00011101011100100101111011011011001000110001010010001011110100010110010011001110011010101011001101011100010001100011100000001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1403[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1403, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000110000010011001011100011110110001111100010000001100111011010011100101011111011000111110110000001101010110010010101111000; 
out1404 = 128'b01011001001001011011001100011101011011111111011110001111001101110111001100000100101110101110110010101011011010111101111000110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1404[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1404, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010111100111010011110000100101100011001100110001100111010111010111100011011101110000010010000101110101001111001010110101000; 
out1405 = 128'b11000010000011101111100101101101100010110011010000000011011100010110011010001110111101110101100101011000100101001101000000111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1405[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1405, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101001011011010010001011010010000101011001111110100101001111001111001011000111011101010110110101010111001100100111001101001; 
out1406 = 128'b00011111110000101101001011101110100101001100110100110001001111100101010101000110011110000011011011111011100110101111011101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1406[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1406, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000100100001001110110100111110100100011100010111101100010101111101000110111001000101111100011101011000001101011100000100000; 
out1407 = 128'b11001001101111011101110100001100011001011000000000001011001111101111111110111001010010101011010010110110011110110011010011001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1407[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1407, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111110000010011111101111001011110111110110101011100101010001010111111000101000011000001110110110110100100110011100011011110; 
out1408 = 128'b11001101001111010000101111110100000010001011010011110100011100101111101010001100110000101011110000100111000011111100100010000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1408[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1408, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011010011101110010001000011101101110001111011111001000010111110001011010011011101101000000100011110101001001111110000011110111; 
out1409 = 128'b00111101001011100111001110011001100001100101001010100100010011011111101000101111001010010011111101000100000100110100110010110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1409[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1409, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111100011101001101101111100100100110000101001110000111101010011011011000111110000110100101100101011100101101001001101100100; 
out1410 = 128'b10010000110110000010001100010111100011111101001001110100100111111010000111011010011001011100110011110000000110010001010110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1410[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1410, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100010001100011000101010100101111011001110101100010110010011101100010010100111111010101111110111100011101110001000111010001; 
out1411 = 128'b01101111000100001100101011000010100100100001111011010010101101101010001101010101010100110110000010101011001101110100010010001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1411[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1411, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000111101011111001011100011001000000000111110001101100101111101100100101101111110001100010011011110110101011111110100011011010; 
out1412 = 128'b11010011100001111010011111010110110111011001100011000000011010111101010110010101011110100000111110101010101000111110011001011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1412[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1412, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010011000100111010001000110100110010101011001101101100000010000111110001110010100111101110010110011010101100000001101011110; 
out1413 = 128'b10000011001101011010111011101010011011100111110101011000010000101100000001110001010110111101001001011101101101111010001000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1413[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1413, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001100100111100011000101010000011000111010100000010101011100110101100000001111011111001111001100111101010001010001010111110; 
out1414 = 128'b01100111101000001011110000010101111011010011101101101100111011000010100101110010111110110001101111000100110001101001100011010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1414[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1414, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110010001001101111000000100100011100100001101110100101110100101101001101100001011100001100000100010110110001001010010110100; 
out1415 = 128'b01101010110011110010101011010100010011110010000000110011010001011001010001110110001011101100100011011010001101011100010111110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1415[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1415, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100100011001011011110111001010001011011101001100101011000010101011010011010010001101001001011101110001110100101101011110110; 
out1416 = 128'b10101010011001011100111111111101110001111010111100011111101011011000011010010110000110101010111110010011011001011000111000011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1416[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1416, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111101100010000010000001110110011100010001001111111110000011100011000000011000011010000101011001000111110000101011000111001; 
out1417 = 128'b10000010101111110110111010010100001101001010011101010111100000010111101100100101010000101111110000100001111010111000100101011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1417[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1417, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100101010010110011110000100001110001110111110010001110011110001011101011101101101001111100010010000000011010100101110101000; 
out1418 = 128'b00000001100000100110010010110010010101011000101100110111001010101101000100110101010001100010100011000011101001000010000011110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1418[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1418, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110100100011011011100010111101111110010010001101110101100010011100111010001111001011100110111101101101010001110100001111000; 
out1419 = 128'b00010110000010011101101000100001000111110011011111000000110010111010101001000010010101101010100010101100001111000111111000010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1419[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1419, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001110011110011101000101101000000100101100000000110000110011010001100011011100100000000101000000000110010101110011010010010; 
out1420 = 128'b00001100101001010100110100110100111111110100110000010000000011000111101111011010000001001100010001111001001101010010101100101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1420[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1420, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111010100000000010001111011111011100010110010101111011011100000001100000111000001011010000000100000110110100010101100101100; 
out1421 = 128'b01101000010001101010000110110101110001111010011000001111001110101001100011001010011011100100011001110101000110011100100001101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1421[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1421, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111000010111000010111000001100100001110000111000110000110010100001111110011111000111101011100100010011111011001110110111001; 
out1422 = 128'b11000011000001000000000101001010100010011111000000111111100111010011111001100100000010010110110101010011010111001011111010100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1422[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1422, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001010110101100100111000011011001110011100011000010000001001010001101011111101000011001100011010110101110011100000111101000; 
out1423 = 128'b10010001100110111010011010110100110010110110101100101000100001010011000100101001000101011101001000111110000111111100111101000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1423[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1423, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001101000011000110100000101111100000110001111001101101111010110011010111000100001101100110010100000100010110110100111100010; 
out1424 = 128'b01000101111011111101011101110000001010101010110001000101101100011110100100001101110100100001000110011000110100111110010011011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1424[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1424, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110000111110010010110100010110011110100111010011011101111110100100010111001111111001011000111010101000010010011110011001100; 
out1425 = 128'b11101011110010000001100111011110101111111001001011010100011100011101001101010011011011110001001110011001110110001001100110000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1425[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1425, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010000110001110101010110111110100010111111010100100010011001011011001000110101000001100010110010110100111100101100010010010; 
out1426 = 128'b10000111101111110001011010011101011111010011000100110100111001000110101110011110001010100000100101010110001011110110111000100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1426[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1426, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101001111000101100100001111110101111000010100001100000111000011111000010010011000110111110101011011100011101000110000001001; 
out1427 = 128'b11101111001001011100110001010100101111100010111110110011011001110100101100101010110000110001010100100111111000111011101110110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1427[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1427, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100010100010000111011100011111000011000101000100110110101001101100111011101101100001010001000110011000010101101001010001110; 
out1428 = 128'b11111110000101011000110110000100111111001000110101111110101001000111010001011010111001000001111010000110111111100010001011101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1428[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1428, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110110010100000100101110011010000000011100011111000110011100001001100110001110001111110011110101011100110100001001110111001; 
out1429 = 128'b11101111011000001110010110110110100000110101110010110111110011000101011010110001010111001000001011010101010001001111011000011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1429[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1429, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010111101001100101010110110000110111010100110110100010000101010110011110000011101011011001011100010100001001001100101010100; 
out1430 = 128'b00010000111100111001001111000011000100111111010000000110001100011111001011111101101100001101100001101101001000010110111011100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1430[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1430, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100010100100110111110111011011000011101110010011000001101111101100011110000111001001001111101110011110100001101011100010011; 
out1431 = 128'b00010101100101010111001001100110001011010011111011111110111010001011111111101101101100101001010000110111010001111011101001101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1431[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1431, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011111000000111001001111010101001001010011101001100100011101110100000101001001110001011101110010110100111000001001000110110000; 
out1432 = 128'b10111000010000111001010101111001010011000111110111100001011111001110100010011011010010110000101001011010111110111001010000010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1432[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1432, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110100111110010000101000000100100001111011111110000110111000000111110100100110011001001100011010010101111011010110011101001; 
out1433 = 128'b10111001001010100001000101011010010101100010011110101110110111011100011110111111000010011111000100010101011110111010000110111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1433[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1433, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110000100000011100000100010111111101110100001011101101110000111001111010110011110111011100010110000011101100110010100011101; 
out1434 = 128'b11010100010100011110100000001000101011011011101010010111111101001010101111010101011110101100101101100101000010111010011111000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1434[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1434, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011110100101111011001101000011111011010110101100100000111000001110100011011011101010011010101111110110110001000101001110111; 
out1435 = 128'b10110101101000001100101111111110101101110110011101101011000000000011100001110110010001111010011000011011100101001101101110111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1435[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1435, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110001100101000011001000111111010111101111001000101111100000001110000101111001011000010100010010101010111110100100110111111; 
out1436 = 128'b01000111101011000001011111101010001000001100101000111011010110010101000101101111001101110100010000110111001111001001110100101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1436[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1436, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011011111001111111001001001110000011100100001011110011001010111110101110110110100011000000111000111011001110110000001011011; 
out1437 = 128'b11101011100001100100011101101001001000000011110001000111001101110110101000010000111010011001111011010110000010111100101110010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1437[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1437, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111111101110100100100000000010010110000010101001101100011110111000010100111011010101110001111011110110000110011111010001101; 
out1438 = 128'b10011111000110000111001111011001010011010110001101001100101101000010010010010001100100101010100011000011111010101011110101010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1438[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1438, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101011111011110111001101000100001111110001101100101111001111111011101110110101011101101000011010100010010011001100111000101; 
out1439 = 128'b11011101001101111010001010010011100100000001010100111101110100001000000010101000011111010001011011110001001010101101011101101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1439[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1439, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110010000001111001011010011110111010011011001000001110010011110010100100110100101001110011111001101001100011000000010010000; 
out1440 = 128'b10001010010101010011100101111011000111010000111111110000100011110010100001011101101111101010011101101111100101001111010110111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1440[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1440, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110100100111100010101001010011111100101011110010111010111001110001100110011111011110000001101001010001100110001111001110100; 
out1441 = 128'b10100011001110100101101000010110001000000011101101101100010011001100000111100111010011001000101110110111100100010111111011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1441[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1441, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110100011111000100000101011001011000011000011000001101111001101001111000100011101010101001111000000001101111011000011100011; 
out1442 = 128'b11011010101111001110000000100001000000100000011101001001100001010100000111011011011000100011111010000101001100110010111110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1442[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1442, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100000110011101111100100010000101110111100000111000111010110100010101101111100000000011011110010011011100011011100111001110; 
out1443 = 128'b11010111101010100110100000010101010110101011010110001010011011100100100011110100011000010101000001000000111010000000100101110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1443[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1443, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100001110001010001001100111000001010110001100100101010101110000010010100000111100101010010111110101110100000010010000110101; 
out1444 = 128'b01101101100001011010110110001111001110101000010000010011110101100110000101101001111110111001110010111111010100001111011110011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1444[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1444, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011111000000011010011111000010001010100100011010110100111111001011001001111111011011101011011010101011111101001011101100111; 
out1445 = 128'b00100101110100010010011010101011011010111011001001010000001010001001001100110111111001000001011010101010010000101101111010011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1445[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1445, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000110100011001001111111100010010011110111000111100100010010101010111110011110101110010011101000011110100010100100011101010; 
out1446 = 128'b01101110101011101011110100001001100101010111101011000000111100010010010111111100100111100110101011101101001000110110101111111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1446[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1446, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101100110011111010010010111101101011011011110011101101101111111110111000101011000100110010110110100110110010011100010101110; 
out1447 = 128'b00100001011011101101111100001011100100011001000011000111101110111111100010010001010011110110100101010010001010101111100101111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1447[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1447, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000011010110100011101011000100000111011011010001110011001100100110101001000011000111001011111000111000000010011011111100010; 
out1448 = 128'b11111010110101100110101010010101110001111111100000001110111000110000101100110011100010000100010111110110010100100100110111011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1448[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1448, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100001110011001000011111010101001100001111010011110000100111010100111000110000111111011000101010111000110111000111100110101; 
out1449 = 128'b00000010011000010101011011001011011011110111101111100010100110000100101110010101000001101101011100101100011110101011001111011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1449[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1449, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111111111011010010011001011000011111100010000010111101001101100001000111011011000010100000000110110010000111111111010010001; 
out1450 = 128'b01001011011011000011000001111100110101101011100100011000001100000101110111010111010000100001011100110111000001110000010010011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1450[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1450, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001001110001111000101111111100001000011111100111011100011011110010111011101010010000111111010111110110100101111110111010111; 
out1451 = 128'b10011001101101000110010010110000111011111100100100010000111110111101011011000000110101100110011110100110101111000110001101101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1451[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1451, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111111110001110010000010011000001110001010000100001011100110100001101000001110111011000110101101011101001111000101101011110; 
out1452 = 128'b01001101011000000000110110011001010101011111011011001011011101101110010101011010110101011100011101111101101001000100011110110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1452[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1452, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100100111011101011101000111001111110001011001011010001011110111001010100010000101111100011001101101011010010011010111001100; 
out1453 = 128'b00110000001000101111011010011111001101110100101110111101100001100011101100011100010011001000111001110100010000101101100110101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1453[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1453, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000010101110010110001000010001110111111101010001001010001101110011010010110001101011100110110101111000001001110100011100011; 
out1454 = 128'b10001111010101101111011100111101011010000111011000001001000001011001111001110111000011001100100100100101001000100011010101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1454[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1454, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011111000111101100101111000010000000011101101000001100000011010001011101111100111011011011111000110110110011110101010001001; 
out1455 = 128'b11110100000001110100000000111100001001011011011000101111111000010010001000011001011001011110101101110111010001111110110110110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1455[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1455, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011010101111000111101101000001110110010110101001001000001110000111101010110110001111100100010110011011000100010011101101000; 
out1456 = 128'b01101101101010000111101100011011000011100101100010011101010111111000101101010100011101001110010001100100001011011010110011010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1456[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1456, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100101101101110011010100001111100001011101000110010110011111100001010000111111100011000111000110010110101101010001010011010; 
out1457 = 128'b10010110110011110100101110100011001110100001001010111010001001110111100011001110010110001010011101001110000110110101010000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1457[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1457, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000110001100111101011101000110000000110111110011100101001110011110100011110000010111000000001110110110111101100100101110111; 
out1458 = 128'b11001000000111111011001100000000101110001110111101010001100110110111000110110000001001011111001010101100101110111110111000010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1458[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1458, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001100100010001110010010001000010110000101111110001000000010010011110101101111110010010001000110111000000001101100010100011; 
out1459 = 128'b10110010110110010110111101000010000110101110000101011001110001101000010110111000101000100111000011011111111001101110100100010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1459[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1459, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111011010011111100001010101000011001110111100101101010010000011010010111011110001100000001100011010100101001011111011000010; 
out1460 = 128'b01011010101001111110111000000101011001111100100011010000100001111000001010010000100101110100000101100010111101110000011101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1460[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1460, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100111010101100101010011011110001101001001111101101011111100101100110100011100000111110101011001100010011010101010110001000; 
out1461 = 128'b10011011110000111111111111111011110110010110010101101011100010101001111010110000001010011100011101100110011011100000000000110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1461[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1461, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111000100110001110010111000001110110101011101010010110110010101111110001000000100011110110100101101101011010100011100101110; 
out1462 = 128'b01101100010100010010011010011111111111000101001100111101000000111111010100110011111001101001010001110101100100001011000010011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1462[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1462, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111101100101101001000110101110101101011010001111001111100010011110011110001011011110010101110101011001010100110100111011100111; 
out1463 = 128'b10111100001001111010101000000000010011000000100000010101010101011100111001101111011010110100010010101111000011111001000001101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1463[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1463, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101001111010111100001111010101110110110111100010111011011101100011000010000110000110101100111101000111000000010111001101000; 
out1464 = 128'b11010011001000011100011101010110010011100011010111100110101101010110100110011001111111110110010011000111110100111000000001001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1464[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1464, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110001100001101101000010000010010111110110100000011000100111100011101000101100001001010110100101000110000000011110010011101; 
out1465 = 128'b10011011010001110000111011000101100011101111110010111000110010100000010100000011001001010001010111001110010001010111010011101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1465[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1465, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110111010101100011111101000011010111001111111011101001101100000010110100111100111111011011011010010101100010010011000011000; 
out1466 = 128'b01101101010101110111101111010010000110100001100001000111011110000101001111100110111011101010110000101111101001001101110100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1466[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1466, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011011010010000100101011000001011110100110100110001000111110001100010101110110110101101001011101101000100101000110001010000; 
out1467 = 128'b11110111001000110001001111011001010101000010001000101000101111100110100010001111110100111010011011110010101111110000101011111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1467[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1467, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011101001011101000110001110001101101101000110000110011010001110011011100011000010101110011000111010000001111000000110111001; 
out1468 = 128'b00101101110101001001011000111000010001110010001011011001011010110101000101110100000000011010011110011110001110101001000100010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1468[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1468, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110101100100101000110000101001111110011010100111010110111110000010111000001100110001100001110100011111001001100010000110001; 
out1469 = 128'b01111000011100010110011100000011111101101100000100100000101110010000010011010100101100101111101011100000101100011111001111010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1469[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1469, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001110011001001011011110011101100100100110011011011000110000100011011010101100101100100000110100111100011010010000100111010; 
out1470 = 128'b11101111110011001100011011101010100100010001100111100011101110111100010101110100110111100101111010110000010011010010000110010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1470[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1470, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111001000100000100100001010111001101011101110111011001110100010110001000101001000010011101010010111101111010000100111000110; 
out1471 = 128'b01101110000100001010100101010111110111110100001011010110101010110011111110100001110100111101100100001001110100100011000011100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1471[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1471, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000000110000011100101100110110000111000111011101111100101001100111011101010010100000001101010101111001100110101110111000111; 
out1472 = 128'b11110101011110010010111011101111000011100111110100111001100101111101011110001001111011111101010001111111111111101011111100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1472[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1472, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011000010101001101011110010101000110111000101011110000000111010111100001011011010101111010101110011100111111110000100010000; 
out1473 = 128'b10001100100001011100011111101000011010111010100100010111110110111100101111101101111010001111111001000101010001100000111100110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1473[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1473, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010110001101001101011011111110001110010001000001001010010100010010010001001011010101001101010101001110100001100000001101010; 
out1474 = 128'b00011001101111011000001001000100000011000011010001110111010000110101011101000011001010110010100010011100010010111100100111001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1474[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1474, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010100011001110001111000100001001010111011101111100100001011011000011011100111111000001010001011001110000111110111111110101; 
out1475 = 128'b00110111101100101100110101101110001001000001101100011111111110011001110010011011110001110100010011000010110110100000011001011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1475[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1475, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011000010001000101111101111001011010010111110110111101111110101010111011111100010111010110100101000101110010001111011100101; 
out1476 = 128'b10011010110110011111101111110010111110100011011001010011001010110001000001010110111011101011111101000100100010000101110010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1476[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1476, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101000100010001101000100101100111010110111010101101110111001000001100010101001011010111010001110100001010111101000010000000; 
out1477 = 128'b00010000001111011011000110000101011010011010011010011101010100010010111001101111001110001011110000111000110110110000001110101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1477[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1477, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101010000010100000010101111111010000001000010100010111001010100100000000001001001011100110010001111000101111110111000010110000; 
out1478 = 128'b10110101100111010011011100100001100101100110101001010010000001011110001101101110110000110010110011110000110111011110011010100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1478[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1478, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010011110001101000000101101001001101011011001011011010001011001101001110000111100101011100000001100001001111000100011111001; 
out1479 = 128'b10011011110010100110100000110100110101010011011011001111100001000101110000101011001100101111101001100001010110010110011110001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1479[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1479, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010111011110100110011010001111111101110100101111110110110010100100110011010011000011001100101111100011101010000001110101110; 
out1480 = 128'b01000000100101000010010100111000111101001110110100101110001001000100001101100100001000001101111011000110010101010001000110000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1480[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1480, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100010110100000000101100010000111110111000001001101000100000000101110111100001101111011100101101011100100101000101111001000010; 
out1481 = 128'b00110101001000110101001011001011101011010000111101011111100010000010111011100100110111101110011100101011000111000001101001001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1481[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1481, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011011011010011101010111111101011110101111010110000010001001000000111011100000001111011001100110010011011001011111111100000; 
out1482 = 128'b01001100011001111000010001101011110100100001011110011110011000111100111110010001000111001001111111110000001101010011000110011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1482[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1482, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011001110101101011001011000111000111101110110000100110000101101101000100110000110000101010110000000010101010101110111010111; 
out1483 = 128'b01101010111100010100011110001011001010011100110000100000110010110100111001100100001000011000100100111000001010010100110111101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1483[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1483, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000111100000110001111000100011110111011111001011110111101000011011001110111011101100011101101111010000110111101001001000111010; 
out1484 = 128'b00010110011010001110010010010000011100000100100010101101101100011110000101000111100011110100000010001011001001011000011001011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1484[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1484, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111000100100010111101101000111001000001000010001010011011011111010010100111111100000010110101100010110100100100010000100011; 
out1485 = 128'b10101110011000101001001101110100011010001000001001011011011011000110101000010100100110100001011100100101100110101100000010100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1485[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1485, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001110010001111010110100110101110011011000010110101110110101011011100001010001101010101100101011011001101111000110001000010; 
out1486 = 128'b01001110101101100101011110000010110110001001000110010000001011001010100110100100101111000100011101100101110110100010100100111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1486[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1486, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110010100110101100111110110010111010000100100111100111101111111111110111000110110100100100101100100100111000111111011010010; 
out1487 = 128'b10111110011001010110011000011111111011101111101000100111001001000001101100001110011100110101110000011000010111100111000100110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1487[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1487, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111101101110111010111100000111000111100001000110010110101111001100010010111110010110000100010111011001111101000101110101010; 
out1488 = 128'b11111110011111100111111011010000101111010111001001000100110001010101101111011001101011110000001101110001101011100001001100110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1488[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1488, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111111111100111000000011100101010001111100001010100100011110010010011000101110110011110010011110001110000011010010001110111; 
out1489 = 128'b10101101101100111000101111110111011011000011100111101101101011111100011100100010110100111010100010100111111010010000001000001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1489[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1489, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010011100001110100100000101000111011111011010000001101010010010101001010001111000001110011111010001110011111100111001111101; 
out1490 = 128'b10001111010000110100010110010110110011000000011000110101001001011110100100110001001011000011101110101101110111011111101000100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1490[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1490, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000011010000100101100111010111111011100110000011111010001100101101110100000001100111001001000000101000100110101100111010101; 
out1491 = 128'b00010010110101101011100100110111111011000101100111001101011110010001110000001110011101001101111001100011011101100100011100110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1491[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1491, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101001001010011010101000011000010101010000111000100000110101110011100011100011111000100000010001110111001101011010101011011; 
out1492 = 128'b01000011000101011100101010001011110010100011010111001100000111011100100000001111111010100110011000010111010010010101100101010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1492[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1492, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111100101001011110111101100100111011001111110010100100001010010010111101010100011010110100011001111100100100010100001010001; 
out1493 = 128'b10000110100001100000001011010010100011111011000011111011000100100101011000111010110100001110000011000111111110010110000110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1493[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1493, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011100000100111011111101111100100101111111000011011011001111001000111111010111110011110001101111100110001011110001110011011; 
out1494 = 128'b00101100111111010000010011011010011001101110001011110110101000100100011110100011010111110110011011110111000101100110100101110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1494[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1494, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000100000011110100000000100101010011011010100010110100000101111110011110011011101110101000100010111100011111111010101100000; 
out1495 = 128'b00111100100010100000100011000110001111010010001000111111101111010100110110001111100101011011101000011010001000001111111001101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1495[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1495, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100001000100010111111010110001101100010011110101001001001111110001110100010110101100010110100100011111101000100111000111011110; 
out1496 = 128'b00101110100010100111000001111101111111111000001110010100011101101011000110001100111011000001010001010110011100011011111111011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1496[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1496, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000110110111110100110001001011110001001111101010110010111010110000011010010010110111101001010100100011001001101101110001111; 
out1497 = 128'b00001101111001000110111011011111110100010111101011111000000100100000000101000011110110111101010111001010100110001011010101101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1497[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1497, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101010101000001101110010000110000000000101111100010111010001100010101000001110011111001011000110100001010000000100110111010; 
out1498 = 128'b00100001101101101001101001100010110010010010111011111011011110100100110011000101101011010101010011101100000011111100101100011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1498[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1498, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100100010001011110111101010001011001101100000001111111000010000101000010100010011110000111100011000001011100010111000010111; 
out1499 = 128'b11000001000111100011001100001100001100101101010100011101000011000110000111001101100011001000011110100000010010001101100010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1499[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1499, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010101101100100000001010001000011010011100110110011001001000010110100001000101110110111100010100100010011111000111011011100; 
out1500 = 128'b00110110101001100111010110010011000001000010011010111001001110101101101011011101111000100011111010000011111000111010100010111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1500[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1500, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100110001111111000011110110000110011101000001100100110101101110100110100000001010111000100100001101101101110011011110010101; 
out1501 = 128'b11111001110001101001101011101000011101010011001101001100001101111010111001011101100000010000111001110000101010010110101000001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1501[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1501, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000111100100011111110100001011000111100100110000010000001100111100111010101101011100110000110001101101100010111001101110100; 
out1502 = 128'b00100101000111111001100110100011001010000010111001100101011010001000111100010011100110001100001000011000100101000011010010000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1502[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1502, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101110110111011001100010011000101011110110110011001010100101100111101110000101101010101001111000100110111000110111100101111; 
out1503 = 128'b11111111101010000010001111111111101010110111100101000000110000000101111100101001011100000000011000111010110100110110010011010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1503[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1503, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101100100001111010001000111000011111001111010001100011001000100000001010110101011101011000010001110001101011000001010001101; 
out1504 = 128'b01101001110101010110011000001100100010000011110100110110010110110100110010001001000000010001010101101110011100010100000001101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1504[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1504, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001110011010111111110011111000011100101110000000101001010100011101010101110110110110110101111101011101011001100101100110010010; 
out1505 = 128'b00101101111001111110111111101001111100010101101001111100110100101010001110000100001010011111010010100100101101101101111111001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1505[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1505, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100001001010100010111111111011000010101100010001010011100101101010001100001001001101000001011100100111100101001011110110101; 
out1506 = 128'b10000111110001101001100101000010011001111000000011101100101010110011110100001001101100111010100010011110010000000100110111100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1506[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1506, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101101001000101010101000011110011101110000111101011100011001011110111010100011001011010110000010111010100101011001000110111010; 
out1507 = 128'b01111100101110110110001001110101111001001110010010110010100100110011000010110101101010100000011100010101110001111000101001101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1507[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1507, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101111101000000011001110010000011011100110111010101011100000000101000111000010010100010111011100100100000111001001111001011; 
out1508 = 128'b01101100001101011101111011111101100011000010100101011100001110010110110010011011010101111001011111001000111101000111010010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1508[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1508, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100101110110000100011110100010111101011010000101100010011001110001000011001001000010010101100010000111111010101000010101101; 
out1509 = 128'b11011101001000101011101101111001101000110101111010100101010100001111000000100100100100110001110000111110001000011101101001000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1509[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1509, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110001001101111010001111110101101010000111011000011110100100010001100110001100001111110000110110101111011111101110111101010; 
out1510 = 128'b00100011100100010000011000001001011011100011101111100110101010101001001001011111001000110110100010000110010100100101110110000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1510[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1510, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010010011011110111000001111000001000010001110001111111110010010110000111101100011010010000001000000110010010010010101111001111; 
out1511 = 128'b00001100111010100111001011100011000101010110101101111111110001101010111010011111101111010000111101101111001110100111011111001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1511[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1511, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101000000111011100100011110111000011000111010100000000001100011110110110011111100000110101111111110010111111001011000001111; 
out1512 = 128'b11010000111001111110101010010110101100100010011000110110111011100101110101100011101001100001110011000000101111100111010001001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1512[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1512, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000101110011000010011110011000111001110001011100011110111110001000001001101011000110011010010000000101011010110000100100001; 
out1513 = 128'b11000011010100001000010110101111100011010000110010110000000001000101111110001110010110111101101110001000101011011001101000001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1513[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1513, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101011111000110011100001111001001000111110001010101110100110011101101111111110110000110110010111100100010101100001101011000110; 
out1514 = 128'b00100001100011010010101100000111111110110100000111001111001100011011111101000100100110011111111000000001000111111000000011111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1514[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1514, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100001101110110100000011110101000111010101000011010110101000011111111110110010111011010001110100101010110010101110011000001; 
out1515 = 128'b10010100001101000100100100010011110111111111000101111000011100100001110110010011101000010010100001000010100001110101001111110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1515[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1515, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011110001011111010000001011100001010100110101110101111111110111010100110101010110101111001100111010111000111000111111110111; 
out1516 = 128'b00110111100010010011011001001101000100111101011010001111110101001011110110111001110000001010011000011111110100001100100000011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1516[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1516, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001011011110010000111100010101110101001001110001001000000011101101000110101101101101011010010101000011111011000101010000000; 
out1517 = 128'b10101011000110001001100100100100001100110000110000001101010000011011111101110111010010000001011101110100101001010101010010101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1517[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1517, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001101110000001111111100011010111010011000011000000011100001011001011100111001101010011100001010010001110010110011111111000; 
out1518 = 128'b11011111100001011111111010110111011010001000101011011101011011100100111110011101110001011101111010110000110100101000000001011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1518[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1518, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100111100001001100101000101100111110011100100011001100101100101000110110011010111101111000111011110011001010111000101100110; 
out1519 = 128'b11111011001101111111011110101101000110100001000110011100000111001001000101010001111001011101001011101100000100100010101110101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1519[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1519, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110010100001101100011111010010111100001000100101001100001111110010001111101011110110000100001001100110011101101000111000100; 
out1520 = 128'b10001100100101000111011110111010101010100001111011000110010111111010110011101000010100001110110111100110000000100001110011010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1520[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1520, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111001001000100100001010101111101010001010111100101110001110001101011011111100001100111111001100000010101000011101100101100; 
out1521 = 128'b01100101000011010011000100011100100011011011111011100000011001100011101000001001111110111101010100111101100110101010110001111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1521[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1521, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011001111100010111010111100011110001110001110011001101010011010100100000110000011101110110110011000010000110101100111110001; 
out1522 = 128'b00001100110111101100010110000110001110001011110001101101110100010110110111110011011010000011111110111001110001000111110100100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1522[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1522, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001110011100111000010001110010011110101000111100101110101011011110100000000001011111011001111100101000111101100101110110000; 
out1523 = 128'b11000101010010011101010001001010110111101101001110000010000010111011001110110100111001001000001110001001110000010110110110111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1523[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1523, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001100111101001010010101111010010001011011111111001100001100110110011110010000100001111100011110110100111110000101001011100; 
out1524 = 128'b00101000011101001101110010110100110110000010001101110110101100101000111001001101101110011001100111110000101101110101011110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1524[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1524, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000101010110011101110110111000110000111011101110011000001000100000111001010110000011001010111000010111011111111000001110011; 
out1525 = 128'b00000000100011111100100100101110001001000010001000110011010100101000111000111111000011111101011110001000000010100110111000001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1525[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1525, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011011111100110011110011110110010100011110100110000001101100100101011101110010010110010011100100010011011000101111111001110; 
out1526 = 128'b00010001111101100100010101001101100110000101110110000101111101100100100110010110000001101101000010101010100101011101101011101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1526[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1526, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010110100010111101100100010011100010100101010011000111010100101001101100111111101110110011101011000011000101111010100100001101; 
out1527 = 128'b11111101100010000110110010000011000000101001100101011110110111010000010100110011100100010010000110011011000100001000100100110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1527[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1527, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011101011111001001011110110011001001010011010101111010010110100001100011010101111000010111000100100001101110111001100000000; 
out1528 = 128'b10100001100001111001101110000010100010110000110100010001110110011010000110001010101111001101001110001101000000110010001111100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1528[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1528, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101001011010111001011101111011111011100110000001110010000100111110010010111010101010111101111011110101010110010111101000110; 
out1529 = 128'b01110011100000100101001111101010111111110100010111000101010110101100111110100101110111100100101100101000101011000101011011100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1529[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1529, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011011010110100001110110010110101001000100100000011011010110101100001101110010100111100001101111010110000110010000000101010; 
out1530 = 128'b11001010001110000010111011111111001000100101110000100001110001011101010100011110101100011111101110001010110010011110011010001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1530[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1530, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000110010101111001010100000000111001000010110100110010111110111100011110010110001110110100110000011011011001010001100101101; 
out1531 = 128'b11001010001001001101111000100111111101100010010110010110011110110101100011011101101010011111101110111001000101010100100010110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1531[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1531, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011100000110010100001000110001010100010010010001010000011000100000111001111101101110101000011111111010011010010100111000100; 
out1532 = 128'b11111111100101101001101011000101100101111010111110001110000000000011111100010000001000000011100110100110001100101111011010010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1532[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1532, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000100001100011001010011101111111110101100010100101111000100100000100111010011010001100111100101111101010100111001111011101100; 
out1533 = 128'b01000001000110111101001011000101010011110011001000000111001010111100111110100011010100001101000010100010101010100000110101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1533[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1533, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011010101111101110001100001100010011111001011110000011010001010011010010000100001100001000000000011100110111100101100011001000; 
out1534 = 128'b11100001001000111011100011111110101110001101100011000110111111001110001100000011101101000101101101011001010011110110010001011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1534[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1534, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001100100010111111100100100011011010011010111001111100000001000110010011010110100110110010011111011110011001001111000110110110; 
out1535 = 128'b11101010110111100100000110001110000101111100011000011111011101100110100101001001010101110110010000011101010001000110010000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1535[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1535, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000110100000110110101001110111001101110011111101000011110111100001011010111010110001111000001111010011110000000001101101100; 
out1536 = 128'b01100010110000010000110111111011000101011010010001110100001101110000001010011001110110001111010100101110111110110011010000000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1536[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1536, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110110101111011000000101001010110000111011001010000011110000010011111001110011011100111011010100100000111001001010000000100; 
out1537 = 128'b10110000000110111011100111100101000010110110111010011000111101011100000000000100001101000110000011111111100101110011110100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1537[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1537, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101100001101001011000010100010101110101000101010010001111101001011101011010011001101010101100111110110001001011001101111101; 
out1538 = 128'b10001010100111000011100100011111110111001100101100111011010100010100010100100010010000010110111101110011110111000100110111100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1538[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1538, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111101001001100101110011000100000100100110001100011110000101011111011010001110110010101011100101111100101001100101011011101111; 
out1539 = 128'b00001111110011000101111001000011001100000011010001100101000001011110001101111110000000100101011000100111111101100111011100000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1539[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1539, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001100111011000011000100111010111001010001001111101110000000011001111001100010111001111000111000110111111111101000010111010011; 
out1540 = 128'b01100001000110010011001010111011001100101010011001000101100001110111100101111110000001111000100001000111011010100011110110101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1540[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1540, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100010110100010110101110011010111101011101100000110010001011100011100000011010001010011110110000010111110010111000100100111; 
out1541 = 128'b10111000010111000111001011001101011110001001110100110100001011110100100110100111010100101010110000011100101100101001111110111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1541[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1541, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111111101111001100100011001010101110100110000010100011010100100111011011001110001101100101110010011110010111011111101001010; 
out1542 = 128'b00101101110110000110110011001000000111011011111011110111000010100100100001001000111011101010101010000100000000101011101100100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1542[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1542, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010101011001010111101110100001011100111111101010010100011101001010001001000101011001001111110010110100111010000110111110110; 
out1543 = 128'b10111011111111101010100111111101111101001111011011100011001100000000100100100011010011110111000110100001111110100101000000010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1543[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1543, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111010100101100011001000001110110000111011010000100010111100010110010110011011001010001110010110111000110100001011111010011; 
out1544 = 128'b01100110010011100110110011000010000010001101111001011111110101010101111010001000101011111111000100101000101100110010101100000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1544[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1544, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110101011001000100010111001111010000001101010001101011100110101000000111111011101100001100011011001011111000000010100111000; 
out1545 = 128'b10100101011101000101000010000100001101111001011100100111000001110101000110010000110100010000000100001010010000110011011001110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1545[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1545, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111000001000100100011001000010101110101100010000000011010001011001110101011100111101001100100110111000100111111001001110110; 
out1546 = 128'b00101110000110001010010010100110011110101101000001010000000011010011011000110110000100101111110100111001010101001110100011111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1546[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1546, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011111111000111010011010101000110001110110001101110000111010100111010010110010100111101011010100000011011001110101111010001; 
out1547 = 128'b10110000000000100101000000101000010101000110010110100011100010101101000000100110000111000111000000000010010110000011111011001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1547[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1547, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101111110100101111111011010000011001101010111111011000111110001101101101100101111011110110110101111001100001010011001010011; 
out1548 = 128'b01010001001001000110110110111001110000000011000010010010010100111100001100110000010110101000001111100000000101010010100111111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1548[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1548, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000101111111001100000010101100100001011111010000011100001001000101001010101100000011010110000011010111010011001010101111011011; 
out1549 = 128'b00101001101100010000111010111010011111011101110001111100111111001001011111001011010110111110101100100110100000110101101100010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1549[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1549, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101001110110100001000011111111000010011001010111001000110011110101101110001110000001110111110111110011100001000000101001101; 
out1550 = 128'b11101011111000110011101011100011010100101011000101100001010000010100100011001100100011100110010011000110001000110100000011101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1550[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1550, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110010001000000101001011111100101001110110110100001111101110101111101011101010010111000111000010110001010111101111100111011; 
out1551 = 128'b01111110000101111101000100101000000100100010110100101001011010110000011101111111110000010111101000000101001101100001010110011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1551[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1551, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000111111101010010110010001111101011001101011100000010000000100001000111010100111001100010011101111100000011111100011101111; 
out1552 = 128'b11110011010111110101000110110100010111110010000011001101110001010100010011111101001110100010011011111001101011111110001101011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1552[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1552, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101010111110110001011001001100010111110100100000111111111001111110101000001110110110000101001100011101001000011110011001100110; 
out1553 = 128'b10101010111101011011001110011010101001100000001100001000100100100010100101101100101011111011001001101001000100011011101010100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1553[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1553, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011110111100111111000010111100001110101010100000000100001101011100111011011101010101111100101110111010110010011101101100001; 
out1554 = 128'b10001010000001101100110100111110111001000100001100000000101101111001011111000010001000010000000110101111101101101000001001010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1554[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1554, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100001100001110010111010001010110111101001111010001001011001100110010101000010000000000110001110100011000111010010101011101; 
out1555 = 128'b10110100110110110001111100010000000000110011110110001000101011100110111000011100101010010001001101111010101011011111001001010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1555[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1555, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100011101101100001101110100001000000010000100001011110111100011101001101101101001110011000000001100000101110000100111111010; 
out1556 = 128'b01101111111101010100010011010001100010001101001111011010000111100011011100000011000001110011001101011100000111110100101010101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1556[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1556, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001111000001011001110000111011001010001110100001011011011011011001101111101001111001101001000111111100001100010000100110010; 
out1557 = 128'b11011110000111011110100111011100110110011010011110011011001011101000001101001001011001101111011001100110001101011101011000001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1557[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1557, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110000001111001011001000110010111001001111001010100111001011110100001110111000001100000011000011000111111001001011011011001; 
out1558 = 128'b00101100011100110110110001101101111001000001101101000000111101010100101100000010110111011000100001101010110001001011101010101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1558[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1558, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100111011110101111010111111010100000101001011010011100110000100011000110000101110010110110111110100011100110001000011111111; 
out1559 = 128'b01111111100010010100100001000010111111110001010001100101010000001100011001010100101101000111100110111000011000100011001000111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1559[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1559, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000110101001100001000011011001100000100100101111110010000100101111111010010000111110110011101101101011000101001110101001100; 
out1560 = 128'b00011101111000100111000101111001001001101100011010011100011000100011110101110000111000111111100111111000101110000100010110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1560[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1560, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100101000101110101000110001011000100011011100010101000000110000101111011001010111111100101011111000100111000000010101000000; 
out1561 = 128'b11110001110000110111100100111001110011111000110101100111001100100001101010111100101100111100111101001011011011100101001010101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1561[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1561, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000010010010110110100000100000001010001111110011011110110110011000111010001010010010111011000110001111000000011101100111111001; 
out1562 = 128'b10101000100010000111000010101101110001000001110011100001111110101100011111110101010011111000100000000001001100001111111000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1562[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1562, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101010101000111001000111010101101001001010000010010001001010100000010000001001000110110001111110011101111011001011010010111; 
out1563 = 128'b10001011001000011101010001101110111110010101110101011011011011101011100011011001110001111101101000010111100101010110100011111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1563[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1563, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101101111010101011111001110100000001011010011100010111011010010001110110001100011110111110001000110001111000100101000100011; 
out1564 = 128'b00110100010100011111010010110000000000000111001001011101111001000110101000011111011000001100110111011111100010010111000001011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1564[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1564, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110011001011111101111101100001001110110100001010101110000110001011000111011110000111011110100111111001010110101011001001011; 
out1565 = 128'b11011110101110111010001011011100000111100011011010000001110101100101100111100111000100001110110010101111101111010010010101001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1565[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1565, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100100011010111010000010000100110010001011101111001101000000011110111111010010100100111001101011100000111001010001101001110; 
out1566 = 128'b10100111110011011000101000110000011000110011010100011110110100011111010001111110111110100110101101011010101100111000010111111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1566[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1566, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110111000101110100111010101110001001111010001011000000001011100100111011011111110011110101111011111011110100110111011100001; 
out1567 = 128'b00000000011000111011000110101011111000100000001100110111010010010111010100011001110011100010101001111010000101010001101100100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1567[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1567, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100100001010101110001000101111101101101111001101001000101111010101100000000100101010101111010011010100111110101001010100111; 
out1568 = 128'b10011001000111000001110010110101001001110011100111111100011101001010111100010101111101111110001110101001011000111000001100101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1568[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1568, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001011110010101100010001101000011010011011110110110110000011111100111110101010011111111011010100110111011010111001111000110; 
out1569 = 128'b10101000001101110100101010111001111000111111111011110001001101011000001101011000011011111000011001011000000111010110001011001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1569[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1569, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110000111001001100110010110001101111010000010110000000001110011111110100100010010101011110010100001000100100100001010011101; 
out1570 = 128'b01011001010000111000001000011110011111001111100001100111001011001100110000110111010010000110110010100110000100111100011000100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1570[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1570, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000010111101101101001010101111110001100110010011100110101110101100111010100011100010111110111111010111110010110010110100011; 
out1571 = 128'b11001011100000101010100010100111011010111111001001010011000001000011011011010111110001100011010010010101110011111110100101101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1571[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1571, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011100110100000100011011100001011111011010100000000000000001111001110111110010000001010011010100101100011111011001001110001; 
out1572 = 128'b00000100111111011110100001001001001000101111010011010011100000111001111110100101001111100110000001100001110110000001110001011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1572[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1572, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111011100100101111101101101101111011100111001000111011011001110001011010011010111110110110001111000100100011100100110010111; 
out1573 = 128'b11011011000101010011010110110110010011000000011010001111001010110000111100100011001111111010011000111010010010011100101011111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1573[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1573, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011110111101010100011001011111110000000011001001110110000110100000100000000101100011011111100110101011110111110101111101110; 
out1574 = 128'b00000000100011110111001001011000111011101001101100010100001010111001101010000001100110000101000110101011011011100010011100100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1574[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1574, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011100101000110011000000100011001100101001011010100110110000001110101111010001100001100011001011011110011010110101111001011; 
out1575 = 128'b11000100100010010000000110000111001111110101010110011011010111011010100011100011100110110101010000100011011110010010100011111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1575[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1575, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010110010001010111110011100101011001100100111111001100001100001010010010110110101111011110011111101111111101110000110111110; 
out1576 = 128'b11100100100001010110010111011101111111110101011100011101010111110001110101111000010100001000011011111101001010100100110111101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1576[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1576, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011000110011100001100101001100111100000001110011010001111111101110100101000010110100011010001100111010011011011011010010101; 
out1577 = 128'b11011110100011100001110101000110100101011011101100110010001110101011100011101100001011100101000010010001011101001010111100011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1577[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1577, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101100101000000011100010010000000000010111101001110010001110111001111110111011101111000010000000000011100000001000100000001; 
out1578 = 128'b00011111101111000111001010111011111101101111010111100010010011001111101100110111011110100011001100100111100101000000111111010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1578[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1578, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011000110111001001101001100110011001110100010001001111011101011100010100011110011111101100101111001111000100011000011101011; 
out1579 = 128'b11110001101100000000010011111101010101110010010000101111010010010110110001111110101000000110001011110101011010110110100001011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1579[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1579, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111110000000100111111110101101010001110111111110010000000111110110001100110100101010010001001001010100110011000010000110011; 
out1580 = 128'b11010111011010111101000011110111001000110010111101101011100011101000000000011011011000100110010000101110000111111010111100111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1580[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1580, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100000010001000001001101011001110110011010100000110101010100010110001010001010001101010100010010100111011011011011100111100; 
out1581 = 128'b00000110010100100010001000111100110011100011001000111000101110011011110101011111001101010111111111101001011101000011101000101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1581[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1581, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100000010101100110000101011100110111101110001000111101100011011111110100101110110000011000111101110010111000101101110011000; 
out1582 = 128'b10010110011101000100110101011010110100000000000101101001001010101011101101101011111000010001000001010000010011001110000000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1582[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1582, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000001011111010100110000111000000110111101100001010110110111001101001100011101110101000010101101011010000100001111000111011; 
out1583 = 128'b00010100111000000101000100101111100100110111011011100001110100110100101001000110100101000001001010110000011111010101001001001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1583[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1583, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001111010011011111000011011101101111001100101011110001010001010100101110010011101111001101111110111001111010011101010010000; 
out1584 = 128'b01110001000010111100011000101110011001101000110100000001101001101011111111010011111110110110111010001010000010011110101010111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1584[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1584, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101101010001111101101100001101011010011010000011011101011001011010010101101010000100110110111010010000001010111101110011100; 
out1585 = 128'b01110101101011010110100010011011010001011000111010000011001100110100111111111101011011101101011101111011001101001001010100100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1585[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1585, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100100000010111101000000110011110001110001001000011011011001101011101010100101110001010100111110011111100000110111001101010; 
out1586 = 128'b10110101110001111110001101011111100100101010001010011111110000100000001000010100000001110000100101011111011001100000110111100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1586[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1586, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100000110111001010110110111110001111010110001101100011010110000111110011011111000111110100100110111101100110001010111110100; 
out1587 = 128'b11101101000001101001110010001101001100111000011011000111110001000110111101010111001101110001110001011100101100100011111001101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1587[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1587, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001011010111000101101011000010100001000001001000000100000001001111110001110100100101001100010111000111010000001000001000110; 
out1588 = 128'b11110010001101000101110001100001011101010011110010111010101001011100011010000110010001101100010000100000101110101000010100000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1588[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1588, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001000010101100000001001100001111011111000100111011100000000010001110110011100010110110000110101010101000010010111110100000; 
out1589 = 128'b11110001000111001000110100010110100100000101001101110000100000011100111111000000111010100101010110111110011111001011000010000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1589[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1589, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001101010111111000011000100101110111001011100110110101001110011110000000010111011000010111100010100100000000110000001100001; 
out1590 = 128'b11110000111110000110110010101100000001100011000111111000110111000110011110011110010010001001011110101000100011011000010111010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1590[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1590, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110100110111110100010100001011010111011010100101100100010111000101000111111010011111011111011110011011101110001001101001111; 
out1591 = 128'b00001010101010001111100000110111001101000000010110001101010101010010000001110110100110000010001000101010100010001110111000001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1591[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1591, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010110011100010001111101101110101110000100101101101110101111001011001101101011000110110110011010111101101110001110110000010; 
out1592 = 128'b01011100101110111011011101010100000100101101111001010010100011011110010011000010101100100010100000110000110001001101011110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1592[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1592, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001000010100100110111111000010011001111001101000000010011100100111111011100011111000100100101110111101110100111001011011000; 
out1593 = 128'b10100101100010000000010001100011101101000010011011111001101001001000100101101100101010111000001111111111010010000101101010101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1593[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1593, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110101010101101100100011011110011100011011100111010011001111001000111111111000011101100000100111001101110100111000011011001; 
out1594 = 128'b00101100110111011000101010001000000001110111000010011100100101101101010000001001111011000101010011010001110010010111100110011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1594[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1594, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011010101000001010011001001101111101001100111100100001110100101011011110010010100000100010111001101000110011110101101000111; 
out1595 = 128'b00011101110111011010010111101101010011001010011001000100101010110111001001111001100001111011101101110011100110100011111111010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1595[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1595, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101101001011000000010111101110011101011010100100000000101111011110010000111100100110100000010111001100111110010100101101110101; 
out1596 = 128'b00111001011000000100101011001111000100110001100101110100110111111000011100010010010111101010110111110111110101010101111011111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1596[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1596, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011101100100101110000101001000001001101100010110111000000000000100000100100110111000111010001011010011001011111101100110001; 
out1597 = 128'b00101011111010101110011111111101101111100110010100010111001111000001110110110011111110000101111000101001110011111010000011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1597[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1597, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011111000010101010111011000111010001000000101100100100101011101111011011101010101000000101100000100110000111111101100011000011; 
out1598 = 128'b11101101001111000001110010001000001010000010010111100000000011110011000111111100000000011100010111110110111100000100100100110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1598[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1598, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101001011010101010111000100100010111110100101001011110001101011011110000100100001001011000011101010100110111111011101000000; 
out1599 = 128'b11111011100011101110001111110001010111101000110110111011011101011010001000010000111110101010101011010000110010010111011011010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1599[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1599, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000001011111111111000000001001100001000101011011101000001100110101100100001001010000110110010101100100010001010101010101110; 
out1600 = 128'b00010001100111010111110110101111000111010110001000011000001101101010010110010110101001111011001110011111101101101101001110110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1600[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1600, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101000101000100000001010111101000110100011101101010001001110001110100100000000010001100010101110101011010011111110010000101; 
out1601 = 128'b00101001001001001111111010110000110000111100101100011000001000110111100101101101100000110001010101000010001110011011011101111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1601[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1601, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000101001110111001010101010010100111110010011111000010011001000001100100101101010111000101110010000001010001100011011011101; 
out1602 = 128'b10110010111000111001000001100110010011011001111011100000100101000000011110100010101110000010010011010010110100111111101110011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1602[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1602, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001100101000110000101011011000111000011001000001101010001011000010110100000110000110011010110011011100011010111111001111010; 
out1603 = 128'b11111011010010111010011011010101010011110000011110110101011011001111000010000100001000111100111111010000100110001111101001101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1603[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1603, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000010000000010100010000110110110001101001001111110011100100000111010111000000111011111100110100100000011000110010100111000; 
out1604 = 128'b01100010010100010010101110101110100010100111010101101000110011001000101010100001111100011011010111001000001110010010101001111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1604[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1604, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100110010000001000011101001110100111110110111101010111001101011011110101101110101000000011000001011101101001001001110010110; 
out1605 = 128'b00101000001101000000111100011101000111010111100001100000101100000101001101001000100011100100000000100001000000100100111001011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1605[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1605, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111000001001110101100001001001101101000010010011110010011111010000101101100010010101101110010111010001000011000000011000011; 
out1606 = 128'b01001010110100001111100110100100001001011000000001110101011000101110000111011001011010011100011100111010101001011111011010011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1606[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1606, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000101000100001010010110000101111110110011101111111101000001111011111110011011011111011101110101110010100011011100010010011; 
out1607 = 128'b11011100011011010100011110011100111101010001010011000100110100010111010011101000000001111000001100101111110010101001101111001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1607[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1607, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010011001110100010011101011000000011001111110010111011001111010101101101000000110001001010001001101000011111001000001010000; 
out1608 = 128'b01011000110110110111011010000111100010010010111010010011101011100100101001010010111101011011101111000001100100001101100111101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1608[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1608, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101001011011100100111110101101101010001110010010010111111010011011001011011000011000000111100000100101100011000111001011110; 
out1609 = 128'b10111110100111000111100101000111001001001001111011100010010101010100001001011001011110110010110110101101111011101001100101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1609[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1609, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011101110100011110101110111101101010011111100101111001110000111101101110010010011100100001100010111011110101010010010100111011; 
out1610 = 128'b00000011111010000100101010111011111001100111101111101001000001110111110100100011011101011001111011110101001100001000111011101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1610[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1610, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001110000000110011110000010000110111101011001111101100110010001101001001011111000110101101110010110111101000100101111000001110; 
out1611 = 128'b10011010111010110001101011001010101001101011100011110110101100011010101010001000001010111111000011011011100111111000110111111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1611[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1611, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100101110010001110010110011101110011000011011000001100001110001111111011101010110111001111100011010100100111101001010011101; 
out1612 = 128'b00001110000011011001011101011011011000111000100111101100101111110101100010000000110110011000010111110111010000000101110011111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1612[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1612, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010100001001111110000101011000010111000000010011000110100100111101110010010000011011101010011001000011111100111101111000000; 
out1613 = 128'b01010101101101111000010001101001000101111110000010111111000011110100001101010110011011110000010111000001010110111000110001010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1613[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1613, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011000111001011101110011110111110110101000000100101110001000100010110111100000110001010010111010000011001101010111110001010; 
out1614 = 128'b01010000001110001011010110000001110010101010010111101100011001001011011000100001001111010010011001110101001110000101100010110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1614[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1614, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110001011010010100110111100011001001000100010101111110011001101110001111101001100010100101000000100000100101011011001000011; 
out1615 = 128'b00110111110011010101011001110000000111011111100000101100001110100001100010001000111010101001111100101011011001010110000101011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1615[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1615, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011011010001001011100011110100110101110101010001011000110101001010001110110111100000000101100111010111110010111000000101001; 
out1616 = 128'b01101110000101101011101101011000110001111100000001111100000011010000110011010100111011010011000110001000011011111100000110001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1616[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1616, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001011100010111010110011001100111111001011011011111000001110010001100110101111100110001010001101101100001101001000110011110010; 
out1617 = 128'b10010000110101111010110000010000100001011010100010011001011101101111111111110010110110001010000111100101000111010000101011110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1617[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1617, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011100111010110111101001000001000101000111110001100011101000010010110011000001000110101000011110101100100000100000111001000; 
out1618 = 128'b11110000111110110000000101001110010110011101011011111110010110111101000100011110110111111111111000010110100010101001011110111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1618[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1618, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110001011111000100000100001111101100000010101100100101101111110000111101100110000100011101000010100000101110100100100010111; 
out1619 = 128'b00010110011101010000010010010000011101100001001000110101110011000101111111010001111001101001111101111101111101100111011000010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1619[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1619, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001100101100111011100011111011110101101001101101000110100011000000110010000001001011010000111011101010011101100011111111000; 
out1620 = 128'b10011100100100111010000001110010000000110110100011111000000010011000010110011110010110001100000001110111000010010101001010011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1620[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1620, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110000010001010110101001011011000010101010110100001110010110111001001100111110000001101110111100101011101101001010110101000; 
out1621 = 128'b10011010000001010100101101100001101110001000001101001111011000010101011101001010000111111010100011100111101000110000111100110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1621[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1621, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101000111000000010001001110100111100010111000100110011100110100001011001100000011111100000111100010111000111101001000110110; 
out1622 = 128'b01100011101110110010110100001011001011101100101101110000101001100011000001011110100110001001010110101000101010000011100011111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1622[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1622, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100010100011100001110100110000000110110011111000000111000101011100111100001011000010010011111111010000101010011100011010000; 
out1623 = 128'b01100101111101010100110111011100100011010111011111110100101101111100100011101000001100010100000001110001110111011100011010101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1623[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1623, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111011101011101011001110101011110110001111010001101011110100110011101111010001001000110011001000100101111111000001111000111; 
out1624 = 128'b01111100111111011110111101010111101010010100001011111000111100101111111010010010001011111001011100001111010101110100110101010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1624[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1624, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100000101110111001100011001111010000110011001011100000101011100101100000100001001001010001001010100001000010110010110010001000; 
out1625 = 128'b01010100110110000111000011111111111110000001001001001101100001010110111001010101100111110010100000111000001110001001101000111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1625[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1625, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011010110111101000111010110000000110111000100101001101111110100100110111000100000001111101010111001011110011111010100101110111; 
out1626 = 128'b10100011010001010111010000011100101110001101000101001110110100111001100111110010101110001011110111100111101101110010101110001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1626[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1626, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000100101000010001010110011000010010100111111001010100110101011110101100010110100011011010011100100001111111111110010001100; 
out1627 = 128'b01100111101100100010100001100011111010010110100001010100111000100101001011001101101111010100011000011110000001001101110100110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1627[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1627, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100101010111001100111111010010001111011100011011110000001011001100011000001101000111101101000000011000101110100100111010111; 
out1628 = 128'b10011110010111001001101101101101011011011001010100111010101011001111110001001101000100100001000001000100000100110010101110011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1628[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1628, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110000010000000011011001111011101001100010101010111000110111110011101101011111001011110111010111101110110111101101111101011; 
out1629 = 128'b11110000110011000110000100001000001100101111001111001011011010001111110110011101011011111010101110000100111100011101001101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1629[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1629, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010101110100100011110010000011000001001010111010100100011010101001110100000010010101010010001000001001011000001111000110001; 
out1630 = 128'b01011011100010111010011001011110000111010110010101100011010011010111001111011110011101010111010001101001001011110011011111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1630[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1630, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100000100100000100001100101001100101100110100010110001110000000101011011111000100010111111101111000101100000111001001000101; 
out1631 = 128'b01001100100010000010010110110000101110011010100100001001000001110100110010000010101010000011101111001001100110111010011101101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1631[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1631, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011111111000000000101000110111011011000000001000000110011000001110100000000011010011110001101100001100001001010101101111011000; 
out1632 = 128'b00101100011000100110010111101011110100111100110110011100100101101011010100100000000111011111111001101100001110010010111101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1632[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1632, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101100011100010100100101010111000101000000001100010000001001010011101111111001010000010010101000100111101011100100111111011; 
out1633 = 128'b01110000111001101011111010111011101110001000111010000010100000100010101000011111101010111001011011000101010011011010100011010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1633[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1633, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101011010001001110111101000010101111000111010111100010100000100011101000111010100010111010010001101010101011011110001000001; 
out1634 = 128'b01011001001010011100101001010111100110001000111010001101100001100111100110001101001111000111110100100010000110101100000011001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1634[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1634, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111011100010101001010000001111001111111100111010010000000000010100101010101010011000001100001011100010111111000000100001000; 
out1635 = 128'b00101001010101011000111010011111001101111001100100000011111111010101110100010110111101010010010010110100011010001110001110111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1635[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1635, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001101010000100010111100010001111000110101010001010101001100110001000110100111110011010111000011010100100001010010001111010; 
out1636 = 128'b11001001100111010000101001001001100010110111000000111001001110010010101100111110001011000101010011001111001011100110001010010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1636[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1636, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101010000110111110111011100100010110111011010011111001101100100001100010100000101011100101000010001110011011001101111001111111; 
out1637 = 128'b01110100101101011010010111110101110110110111101011011000111000001001101111111010000111000100010110101111101100101011010000001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1637[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1637, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100001111101101010011010010001000010111001011101100100010011111111110111001011001100100011101101010110111000001011000111000; 
out1638 = 128'b10100001000000110101011001000010000101001011110010011001100001110101000000110011101010111011111000110001001101001110011010100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1638[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1638, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010111111010100010000000101100011100100110101011001010100010101100100110100100011000001001011011010111101001101001100100110; 
out1639 = 128'b00111111110010001101000000001100010000101101100100000000001101000100011010111010110110100001000001000011100001111100110100011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1639[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1639, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111100100110001101111100000001010000011101011111011100011011001110001000100001010001101110101110101110111000000010000000100; 
out1640 = 128'b10111111010010001111001011010100001000000010111101100011001111010100011000000111100000011000000011100110101111000100100001100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1640[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1640, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001100010101011011011010110101111010000011100001110010111010101010110101110000011001110110110001101111010010110100011101000010; 
out1641 = 128'b00001000010000110110100000110010110111000100110000000110001110100101011000010000100101010010101101100111011011011101101000111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1641[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1641, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100001001011001010000111001100111100100101100010101101101000010001110011100100001010001110111100111100010110011010110010111; 
out1642 = 128'b01000011111011010010011001000101000011101110100001010100010000000001110010110000000100101110001001001110000110001110110111101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1642[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1642, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000001000000101111110001101100001011011011110011110001010111100111000111111111001111100101010001100010111111010101111000111; 
out1643 = 128'b11101000011000001001110011010100001110010011100100101101111100100001100100110011001001000111001010010011011000001101111000000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1643[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1643, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100010101011010111011110001100010101011001011010110000100110010010110010011000111010111100111010110011001001110000000111010; 
out1644 = 128'b11101001000010100000101010001011110001100100001111000101111000000010100111010111110100000110010000010001100111000101010000010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1644[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1644, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110000000010101001010000001001011101000101100000000100001010010011110111010111010111011011101111010100101001100110011010110; 
out1645 = 128'b00111101001100110111110001011001100001001111111001010000111001101111010000000001010100011001111011111011011101001100110100111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1645[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1645, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011000100001101000101000001100001111000011011000110101111111101011000011000111000011111101110101000001011101110101111001001; 
out1646 = 128'b11000111101111001010111100011111000101100000110100101111001110110110001001111111111000101100001110010111010111101100110100001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1646[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1646, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100011011011011101110100011010100001011100100101110000011000000100111000011111111010001000100111010101010011010001001100000; 
out1647 = 128'b11101100110010010100000111110010011011110110101110111101110111100111101001011101101001101101100110010010100010111101000011011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1647[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1647, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000111000110110110110001001100000101001010100101111100001100001100010010001101100011001111011000000001101100001001111001100; 
out1648 = 128'b11000001101101101011011001111010100100111000010000011101001001000111111011110111010100011111100111111010111001100100100010000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1648[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1648, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011000111111101011010111110100000111001111001011010010100101110111111100001100110111101111111011100011000010110100011010000; 
out1649 = 128'b01010011110011110100010111000100100110111000100100011010010010001110010110000010000001001001000011101101001101000101100000101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1649[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1649, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111111000010011110110011101011001000001010101001000101111011101011101000101001100010000001001010100000011001100110100001001; 
out1650 = 128'b00100010010101011001000000110000111111111100100011100110010001001011010011111010100100111000001111101100010000001101000101010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1650[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1650, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100001011011101001100000110010011100101011000001111110001001100010100011000111011110010000010100001110110110101111000100010; 
out1651 = 128'b11101101110101001110111110001111110110000000100101110000001011010001101001100100000001011101000001101010101100100001010100101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1651[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1651, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100010110001111001011001110101111101001100111000011011101111001001111000000001000111001000100100111100010011001101000010011; 
out1652 = 128'b10110010110101001110001101010011101011000000001110101000000110111001011101101001000100111101000111111000010111101001111000011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1652[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1652, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100011000000010110111000011101010001001100111001101000111011010101010100100010111000111010011011110011100011001000100111010001; 
out1653 = 128'b01101011001100110100101010010010000100110111000111001110111000000011111100100111101110101010010000000110001110000000000000101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1653[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1653, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001011110100100100101111101001100111111111011010110111111011011001010011010100110000111010100111011100110001111111010110011; 
out1654 = 128'b00001101100100111110111010000100001101110101000010001000110010011110000011000101100010011111011011101000111000111110110001001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1654[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1654, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001010111101100000000010000011100010111011101101001011111110000001110000010010010110101101001000001000111010111101010010000; 
out1655 = 128'b00000110100001010100000110001100110110010110001001111101101000001111101100110011101100001101010011110111100110101101001111011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1655[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1655, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001111000001010001110100000001011000100111010000011101100100000001100000010001011100011001101001011110000100111111101101100; 
out1656 = 128'b10101111001101110101111111111110010111011101101111000011101011110110100111110111011001000000010100011001100111101001011100010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1656[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1656, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110100010011101110011000100110001000100101000100100100010110011110010000110101100000100101011100010101010001110000000101010; 
out1657 = 128'b10011010010000101011000001000010101110110101010000100110100011000000001000000001000111001100011100000011011000100110010011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1657[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1657, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001101010010110111110010101111000110010000001110100000101001101000010010101100110100010101010100011001010001111110110000000; 
out1658 = 128'b10110111000010000100111101100100000110011111011110100011001111111001101001100010111001000000100111101100001000010100010110000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1658[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1658, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000101000100110111000100001001101111100101010000111111011110010000011100000111100011010001000101111001000010100000000100101; 
out1659 = 128'b10001001000101101011110000111011100011101010010001100101100010011000010010010000101001001010011111000100111100000001010110111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1659[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1659, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111101011011110100110111000000101101110000110010110101111010001010101111010110111110000011110011101110010010011010110101011; 
out1660 = 128'b00001010010101110100000100010001000110111111111110110100100100101001011100100101011111010101111010011111001000010001110111001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1660[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1660, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101110001100011000110100001001101101000000011000001010001001010100100000101110000101101111000110110000010111001111010111001; 
out1661 = 128'b01100000100110111101011000110001111010010010001110000011110010011100011000111101011100100000011101000001110101110101110010011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1661[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1661, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010010001001111000100110000000000110100101110110001000000100100001001000111101011000110011110001110101100110110000000010010; 
out1662 = 128'b11000000100001110110100100000000100001100010111101010111000001110010010000100000001011011100111100001101110100000010111111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1662[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1662, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110011111110001000100111101010001111101100010101110101101101100100000010110111001011100010011000010110011111010100111000000110; 
out1663 = 128'b11100111011010000000011001001100010011001011110111001001001000100100011010000010101101011100000100111100010101101010011010110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1663[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1663, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110111110101000011000101110100001110011101101110000010000110111110011000011101011000001010000100000011001011000001100000100; 
out1664 = 128'b01101111110011001110111100111011011001101111100001110011010101111000000010110100001110111101000100111100010010111001011111101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1664[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1664, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101001110100001111111001010101000100000111100110010110000101000100011100011110110000001101001010001101001110011111010001110; 
out1665 = 128'b01100100110101011110000010101011101100111110111000000001111010101010001011101011000010100110010101100110000010100010100100101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1665[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1665, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001111001001100110000101100101101001011011011111110011001000110111100110011111010101001111101011110000001000011000000101010110; 
out1666 = 128'b00000001100101001100001001010001010101111011110001110001110101100010100000000101110010001001101110101001001011101100011010001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1666[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1666, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110100010110000101100010001101011011110000100110010011000001100010000110001110111001010000111000100000110101100100111000100; 
out1667 = 128'b11110100100110001101000100000100011110010110000011010110101010101100111010111110010001101111100111010110000110010001011111100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1667[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1667, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111010001110001110101010100011111010010001110101000001011101100101010100011100010110000010001010001011011110001010001011100; 
out1668 = 128'b01011001010011101001101000001010100100111110111000100001010011000001101000000111101110100010000110111001110100001100110000001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1668[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1668, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101001101001111011000000010001010001100101101000000110000110110100000110111000000010110111010110111100010000010001000110001; 
out1669 = 128'b01111100001100011001111100000011101111111110100010000110001000010111010011000000000101111110100110000001011000000101000101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1669[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1669, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000011111000000001100010001101010001011110111110110101010010010110010100010011001011010011111000001001010000011100101010100; 
out1670 = 128'b11111100110011001110111110010010100001110101110110010001100001101100111010011100111010010010111011000101010001000101101111110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1670[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1670, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010000000100011110001000101111011010111001010111011111100111001100110101111111111011111101001001010010000000100111111011010; 
out1671 = 128'b01100000011001100110000000100110000111011110101111110100101010010011101101001000101011110000011011001100110010101100010101010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1671[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1671, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100000000111111010010011001011000101111100010110011101110100111101010011100100110101010011001101100111100011110010010011100; 
out1672 = 128'b00110101110111101010010100101101000001001100111110101001001110100011111000111011101011110000100100100010101001111100000101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1672[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1672, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111000000000111111100111111001101110101001110011100101100010011000100010100100110111010001111110000011100110011111101000101001; 
out1673 = 128'b10001011100110101001111000101101000000001001100110010001011001101011001001000111111100110100010011011101001110100100110010000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1673[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1673, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001000001101111101000100010100100110011100101011010000110101101001000001100101101110111010011001100000000110000100010011110; 
out1674 = 128'b11110101111000101100101110101000011000110100101011110100111010010011001001101011100000110011111010110001110001101111100101110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1674[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1674, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100111101111011011101011001101011101110100101001100001010000111011001000010111010100010011110101100100010100101101111001011; 
out1675 = 128'b10101011110011011111001111101011010011101011000111110011010000101000111101011101101000111110010111010011000110110100001011100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1675[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1675, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101000011000110100010111000000011101011110100101011001000010100011010011000110010111000011000101010001001101011011001001111; 
out1676 = 128'b11011100010010111011001000111111101111110000011111011100000111000011101100011111000100001011110110101000100110110011011101001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1676[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1676, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100100011000001010110101000011010110001011100000101100011100110100110001110010001110011010011010110001101011001011111000000; 
out1677 = 128'b01010100101010100110011010110000000111000101100000111110100111111111011011101000001000011110001010001010100010000111110110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1677[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1677, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011000011010011111111011011101000100100111110110100011111011110100011110011100011111000111000010110110011010010010101000101; 
out1678 = 128'b10111010110111000011000001010011011110001100101011010010001110110100110010111010000001111111100101011101010110101100011111001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1678[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1678, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101011101000000110111000000111011000000011011001101101001001100100011010011000000110110111101100010010101001110100010011011; 
out1679 = 128'b00001101011101010001011110001100001000011010000110110010101100011001001111000011011101100110001010011111110001011011101111000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1679[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1679, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001011001001001100001000010111101101000100110110100100100111001011011101111101100110010110001000011110001011100110001110001; 
out1680 = 128'b00011001110000010101010010001110000011000101100100100100010001111000110100001011000101011001010000000111010110110100100111010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1680[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1680, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001011111101111010101110010110011111010011101110111010101001111010001000001011010001110011100010000011000000101100101010011; 
out1681 = 128'b11100011111011100110101001010110011111101111000100000101001101010100100000000101000011110100000010101101111010010111101101111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1681[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1681, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100010000010111111010010110011100110110000110110100111001110100110000011000101001101010101001100001010010000110010011011010; 
out1682 = 128'b10111010000011110010001111010100011000000100100011101111110110110000010001000101110011111011011011011001101110011100001100111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1682[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1682, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110011001000010001010101000011001010111001111110000110110100101100111101101011010101101011000111011011001111010001011010101; 
out1683 = 128'b11011011000111101011100111101111010000000001010011010000011010111101010110000111110000110011101001111100101001101100011010011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1683[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1683, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110111110001100000111111000111110000111000101111101100100100100101000101111001100111110001110011010110101101000110100011001; 
out1684 = 128'b10011010010010001110001011101111110001100001101111011111001000001011011010100000011000001000111010010001001001000011111111011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1684[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1684, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000011110101001101111111110111100111001111001001010110010010001100010001000000100001001100011001001010000011100011110001011; 
out1685 = 128'b11110011101111110001101101011101010101111001011111011101111110000101010010100010111011100010010001010110101100100111100001001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1685[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1685, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000111011011101100100111011011110001101001001100011100000100000001000101010100001110000001010011101010011000011000001110010; 
out1686 = 128'b10101111110111100011101000101101011001001010010000110101111010010000111100001100101010111101010001010001111100111101100010100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1686[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1686, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101000111001010010101010110110001001000010111010111111000010110000001111011110100010110110011100101110101100010101101100010; 
out1687 = 128'b01001101011011000000011001100011110010100010010000100111011100111101100011000100011101010100110011010000000111001101011110100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1687[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1687, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000001001110011011011100111010101000100100010011000011101100100000000000000111010010111110111101011001001100011110011001011; 
out1688 = 128'b00010011001110000110000110100100000111100000101000000101101111110000011001110001011011001001110010111010110110111101111000101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1688[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1688, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011000110001100100011111100010110100111010001110001000010100100010010111011010101100001111100111101101111000110110100000110; 
out1689 = 128'b10110111000111110100010110101010100101111101110111011011000100101110001110010000000001001111101110110110010010000011111100100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1689[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1689, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101011101010111000100111110110101100000010111100100000100001110111000111010101111110011101100101100001001100000101001111011; 
out1690 = 128'b10001011110000110011100011110000011110101011101110000101100111101110011110001111001110001001110111000010111101000010011111000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1690[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1690, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100101110010001001111001010000010101011101001110011110101100010010011101110010100000011111010111011010111001110010100010100; 
out1691 = 128'b11011010111110111101000111101111010100110110111001101000011100001111001111110110010001001001000000001001011000100000100010101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1691[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1691, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011001011000001011101010111100010011001110001101111110011111010111010110101101110110110000110111111011101111110100001010111; 
out1692 = 128'b01011011011111010001001011111110010010100000010110000101011101000001111010001101101110101010110001000001010100000001100001011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1692[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1692, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101110011101111001110011111001110001111101010011100110101111100110111111101100110011110000101110011001111010111111100111111; 
out1693 = 128'b10110101000000010101101100111110101011010001001111010001101111001001100110101001011110101000011000100110011100111010010001100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1693[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1693, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011011011110110010110001111111011011001100100000000100010000101001101110011111010101110000110101111101110011110011111100000; 
out1694 = 128'b11001111000100011010000111110011000001101001100100101010101011000111101010100001010000000001110011000101000010000010100010110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1694[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1694, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010101001110111100101100100111110101010111100100110101000000010111011011000011000010000011101111011111000010011010000110110; 
out1695 = 128'b00001001011100001011010011001011010011001011111100100111010000101000011000010110011101101010000111011010011000000010111010110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1695[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1695, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011010001011100111100011110000010010010010001000001010011000001010010101110011010001100101010110010000111011111101011101010111; 
out1696 = 128'b00111001101010110011001101101011001111100011001001110010010000111101110111110101110100110000011000010001010111001011001001010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1696[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1696, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001100000110100011110001111000001111000000111011001010011110011011010011011100110101001111100001000110010001001101000101000; 
out1697 = 128'b00110000101100000110000011000101111010101011101011101111110111011111010011000011101101111101000001000111110001110011111101111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1697[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1697, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010110001000110010000001011001010111010000001101110110100101000110100111100110100101111001110110100011010011100110010101110; 
out1698 = 128'b11000000001111110111001000111111010000001100100000101111011011110101000000101001101010100101110010011000001110001111011100101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1698[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1698, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100110010111000110000010110111011001111100000100101101000111100011100011111100001101000101111011111001011010000010011001000; 
out1699 = 128'b01111001100010110011101101100101110111001000000101110110111010111111001100001010010010100100011110001000100011111101110100100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1699[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1699, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110001001000001000010100011110100001011101111100101111011111111010110010001100100001000011010101010011111011100101001110101; 
out1700 = 128'b01001101110101100111001100000000010010000001010010001111011110111011111010001100010110111110110001000101110100100001111001111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1700[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1700, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100001101010001100110111010110001000011000000100101111010100111110000011111011100100110000101101000111101111010100100011110100; 
out1701 = 128'b10111011010011101011110111110100101011100000110011010111010010001101000100001011110010100011001000111000101100011010010011010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1701[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1701, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011111010101000100111000100101001011100000100011000011110010010010011010111100001000111101000101001011010110011101000101010101; 
out1702 = 128'b00000101001011101111011001000011011011000110010011001111111100110100010110101101010111001001100110000100101101000011011101111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1702[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1702, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100001000011101100000001001111100000101111100100001111001111000010111111100101101101010101111110101111001111110100011110111; 
out1703 = 128'b10011111110011110001001010001001010001011010000111110010110110100100001111100111111110100100100011100100111001011011011111010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1703[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1703, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111000111101011010111111010000101010111111001000001010010101100101110001100110010010100100100001101001111010110100110101100; 
out1704 = 128'b11111011010011100001100110011100101000000101011101110001010011011110000010010111011111000000011011001101010111011101011110101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1704[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1704, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000011011000110100001001111000011101001101010100101000001011110001011001100010001000010001100100001000001100111111001011010; 
out1705 = 128'b00010100001101010110101000110010110101000001011100010011010111100111000101000011111000111101110011111000001011101011100001110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1705[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1705, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000101011101010111010111111111011111111111100100101110111001000000100101001111000110001011100011101101010110100010111100110; 
out1706 = 128'b01111111111110100000000110100100000101101100010010110001000100011010011011110011000010111001001010101001001011001001001101010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1706[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1706, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100010000101011010010111011010000000010110011100100101010100100110010100100011101110011001110100110110110010100110011010111; 
out1707 = 128'b11010001110101011010111100000001110100010101000010001111111000011100001101100001110101101101111011011001100011101010001010001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1707[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1707, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010000111001011001110011111001010000101001101011011111111010000111011110000110001111000001110000010000100001110010000010110; 
out1708 = 128'b01010010001111111000100010011001000100010010100010101100000111101111110100111011010000101010101101010010000110011111001000100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1708[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1708, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110110101101010111111010110100100110011010000111010011001111101011111000010011101011010001110010101000110110000100001000111; 
out1709 = 128'b00001011110010011001010111000100000100001010010100010111101011011001010110101000010110000001001011100111111101110011010010100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1709[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1709, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110010111011110110101000000101110100110101101110101101001011101011001110101110100001100010100111110111110001100011100111111; 
out1710 = 128'b00111010011110010001110110110010001110000001011011011111101011001010000101001001111010111010010101011101000100111110100100010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1710[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1710, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100100100100101111000101100110110011010000000001100011011000000001110011100011001110101111110111101000000000110111110100100; 
out1711 = 128'b10011010000010100011010101111000110111111010111000110010010100111110100111000000101111110011001101111010110001010000110001111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1711[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1711, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011010000111011100101111110010000111110101110110100100110111010010110001101100011110111011101110000010110100010100100111101; 
out1712 = 128'b11110101000011110000011101100010010011100000001110100100001001010110000001000000100010001100111100101000110000111010101010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1712[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1712, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001011010111101000011101001010001001011101011110011111000100011110110110110011110011001111100000010100111101110000011011111; 
out1713 = 128'b11011000111100101010010001100101010101001111011011010101101001010011110011101001111101111000000010110101111011100100111011011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1713[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1713, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100100000010011001000011000000010010111111000101101111001100010111111000011111000111001001010100010110000000011000000111000; 
out1714 = 128'b00110011101110100110110010100101000101110100001010111001001010010111100011111010111111011000100011100010101001000000100100010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1714[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1714, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001011100111111101110101100010100101010101110011010101010111101010011011011011101001101111001001011100110110000010000111101; 
out1715 = 128'b00101100001010000000011101111111010011000001011111100010101101000111101110111001001011010000100101110111100111010110010000001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1715[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1715, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011111000000000101111000001010101011101011110010011011110110111010100001100111100001100011110000000001011101001111000100010; 
out1716 = 128'b00110011011011100101000000011111010101101011010101011101000001110101010100000110011011001010010101111100111011000100101000110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1716[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1716, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011100111000011110100100010110110111111000001001110110110110100110011001101111000000110010110110001000010100100111000100011011; 
out1717 = 128'b10000111010101010110100000000111101011011100000000010100110000001011100011101100110001011001111011100100001010111001100101101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1717[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1717, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011110101100000101000110111011011101101011011010111011110110100001110010111011011111111101110100000110100101110011010010100; 
out1718 = 128'b01101101010101001001011110100011001000110000010011011100001100101111001001010110001110011111100000000111111100000110000101010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1718[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1718, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111000010111111011110110000111010111010111110110001010100100001100100110110100101100110101111110101111001101101111101000001011; 
out1719 = 128'b10111011000111010010001101010000000000110010100010010011100101011011100011010000000110100101111111100101101110110001000001010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1719[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1719, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100011100010110010010111110011110001110001011111011010100111001000010100111110010010001110000000011100101001011101100011010; 
out1720 = 128'b11110111011100100100011111111101011001011101100111000111001101000010100100001010100011100110011011101100000111000001101100010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1720[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1720, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111000010000001011111100111011011011111101010111101101001000111111001100111100011000110101101010001111000100100110000100110; 
out1721 = 128'b01010100011001000100101100101011101100011000001010101101100111011010000000111010000010001101000001000100001101101011100010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1721[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1721, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001101001101000001001000011101111010011111010000100101011001001010011000001011000101010011011101101111110100101110010010000; 
out1722 = 128'b11101000010101011101110110000000111010101100010010110001101111011111111001011110110010010001101001000101000101100110001000111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1722[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1722, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011010000110000101101011101100001101010011110110011010111001100011111110000111010010101001100000101111000010110110110001100; 
out1723 = 128'b01011111010100110001110110111100001000011111111101101000001000000011010101111000101101000010010110011011101010000010110001101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1723[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1723, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011011101010111001000110000100110000001111001011111101011111010011000000010000001100100001111010001010001111110001001111011; 
out1724 = 128'b01101101010110001100001011111101101011001110100010100110101111110110000111100000011100001010011010100101101001000000011110000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1724[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1724, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111011110011001001101011011001101111001010000001010100011111111110010100011011100110111010101111001111100001001110100000100; 
out1725 = 128'b00011100110110001110100011110110010110100111001010101000010100010010011111110000010100000110000110010001101110010111101001111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1725[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1725, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001000000011000001010100011010101011000110110011101110000101011101011101010001001100001101011000111011010000000100100010110; 
out1726 = 128'b10100110101010011000101110000101101110000100110011100001010000000100101110001000100100000111101101100100111101100110110101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1726[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1726, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110100110001111011111010111111110000110111110000111010001010110110000011100111111010111000010110010101001000110101101111101; 
out1727 = 128'b11010011100011000101011111001101000110000011111101001110001111101010111001110000011101111100111000100000001111110001001000000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1727[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1727, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010101100101100111111001010011011010010111110010001100111100010100111000011101001110111010100110010100001111011011101110001; 
out1728 = 128'b01001101000111011111010111010001010001010010010110010101011101111010101000110100011101100110111001000100010101011010011101011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1728[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1728, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111100010100110000111010111101010001111010010000100011111000111111011100010001011111001011011001000011011101010111100000011; 
out1729 = 128'b10000010111011000011100101011101101111001110110010101010010011011110001111111100010000101010011110011110011001001110100111010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1729[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1729, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001011111101000000001000010000111110111011010000011010011100111000001110011101011011000101001011010110011010011010011111111; 
out1730 = 128'b01110010111001000010011100010100110010001011100101110100111001001110111011001101100100110000011110000010101111101110011101001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1730[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1730, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000100011101001010000110010000111010111111111010101000111110100100110101100011111000010101011110110110000010001011000111111; 
out1731 = 128'b10111010000110110010011101000101100000100000101110010111000111000100110111000011010010111001100011011001001101101001101110110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1731[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1731, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010110010001100001010010111011011001111111101110111100011100110110100000111100010111110001111011000110100100111100101100111; 
out1732 = 128'b11011111111110010101110000110111011100111010111010100101001110011100100100101101010110000100010001111101001111001011010101111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1732[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1732, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110000101010110101010001010100110101011111101010101011011000110100101100110101100000001011001100100101100010101110001011110; 
out1733 = 128'b10101000110010001101111011010010001000001000101110010011000111001001111100011010110010000010101011001111011000000101101001101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1733[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1733, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100000110000010111000001110010000011001000010101001100011110110100010110001110000110000100101001001110010010100010010001010; 
out1734 = 128'b00011110101000100010101001110010111000001100110011100111100001001011001010100010011001101000001001000101100011111101011001001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1734[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1734, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111101000011111100010101010111101001010101010111011100100001011001110101110111000011111101001000010010101011000111101100010; 
out1735 = 128'b11000010100111101000000001101001101110001111101001100011101010010111111111010101001010001111101010010100011101011011010100110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1735[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1735, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100100011110100010000101000011111011111001000000000001000111100000000111101110001111000001111011000110111000110100111001111; 
out1736 = 128'b10011100001111111011110001011001011111100010100011111101000001110111100001110110001001011010001001011101011100011010001011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1736[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1736, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101100011010010001011101101100100100110101000000111011011000001101001010101111011010100110010011100110000011101100011010100; 
out1737 = 128'b10010111001110000010110100100000101100111110010111110111100100001111101001100001100011010111100101101000001000011101010100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1737[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1737, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011001110100011111010011010000110010000000110000001011010100101111010010011000011001000010011101000011011001001110001000101; 
out1738 = 128'b10100010010010001011111010001010100100010100001110111010111110011111101011101001001011010110110100110011101110100111000110000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1738[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1738, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110010110111001011011101011111001000101010011001110101010110111101001110000101110101001110101000101110000100111110111000011; 
out1739 = 128'b00100000110101000000100010011100101110111000111111001100110001011010011100101111101111001110001111100110110111011110101000110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1739[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1739, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111101011111000100101010101010000011011101010000111100000100011001110110110100000100101000111000110001111110011000111001011; 
out1740 = 128'b10000000011011001000000100011111000110101011001100011011000000110110110000110000111100011110101000001001011001000011000101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1740[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1740, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101110011101110010100110101000101011001001000110110110011111011010110100001110000010100010000110110001111111100010110011001; 
out1741 = 128'b11100101101110101100011011100000111011100001011100010010110100100110010000001010100011000110110001101011001000111101011001100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1741[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1741, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001011011110011110000100000001010001011001011001010111001001110000001011000000101000111110111010000001001011001001111110111; 
out1742 = 128'b01001110111110000001010111110100110010100011100100111110011101011100111010100001101010000001000000011101011011000100110011011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1742[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1742, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101101011001011001010010110000001110010000110000111101110000100110000101000100100111011010111110000010100011010000101011010; 
out1743 = 128'b01111100100010100011111001001110101010110011011101111001000110111110010001111010010111100110101111001000010000001101111111110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1743[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1743, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100011000000010011001100000000010001011000010010100010101011010011000001010000010100010001011000101000100110111011011000010; 
out1744 = 128'b11101001100000011001011111111011001000010000101110001111110010101111010010100000110101100111101111010001110100110011001110000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1744[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1744, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100011100101100000001011101100100000110011000101010000100100010110101110010100011001011001110110000100111010101011010100101; 
out1745 = 128'b10011010000000010100010011011000101010110111010111000111100011001000111101111111000101100111001011101011011100001000001110100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1745[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1745, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010010011110001010010101011111010100011000000101000100000000010011011110001101101010000100001100111000110010010001111000101111; 
out1746 = 128'b11101010101101001101111110111100011111001101110010011001100001110110100110101000010000000111000101000111001101000111101010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1746[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1746, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101111000011000001001111111111100010011010000011110100001110010011100000100011100111100000110010111101110011010101111111110; 
out1747 = 128'b11011010011001011111000111011101001000000001101010111111010100001000000000011001110100000011111111111001110110110001101001010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1747[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1747, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111010001001110010111011011001001001001110001101000000101011101100000101010100001110000010101000011100011100110001010010000; 
out1748 = 128'b11111000001000000101110010011010100110011010011000100110001110010100101010010011001011101001111001001011110001111100111101011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1748[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1748, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101101011010111010110110001000111001010110100010101101010100101011000101011011000100011110011101001000000100000110001000011; 
out1749 = 128'b10110000110001011110100000001110010100101101110011111011100110010100100011000111110011001100011101001010100111000000111110011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1749[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1749, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000110000000011001011111011111100111110011011110011101001110000111101101010111011110111011011000011011111000001110110100000; 
out1750 = 128'b11010001111011111001000001011000111110001110000110110111110001110101000011111001101000101010000011111110010010110100001111111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1750[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1750, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110011011001001011010111010000001100101001101110110001101110101011100111001111101110000111011001111110110001000000111101000; 
out1751 = 128'b11110100101101001011100110111000001110101000101110011001110011100001000100111000010111100100100000100100010110000111010101101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1751[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1751, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000111001111000010111010100100000100100011000000000110111111000001111001011110110011011101011100001101101101110011001110110; 
out1752 = 128'b01101100011001011110010110010001010010110011011000010100111101000001010011111111110101000010000001010100010010001000100010101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1752[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1752, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000000111001100111000101011001011011110001010111000110001100110000010110000100100110001010110110001100010001110110111001011011; 
out1753 = 128'b11011111011001000010011101111011001100010010111010111000011011110000010110001110000101110101110101010100011000011100101100110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1753[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1753, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000011111110100010111101010010011111011010101010010011111101011100110000111110101110000000010110101110001010000001100001001011; 
out1754 = 128'b01100111111101100010001110101100100101100111011011011011001110110000011101010101001110111011100001001000111011000111011110101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1754[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1754, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110110011001110100010101011010011111110101100101100110001000000011001011011010101011110111101101010110010110110011000100001; 
out1755 = 128'b00000000110000111010000001111101100111110111101011010000011010101111000111000110011011001101101001001011101100001111000011110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1755[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1755, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010001101001100011011110110100110011101101111000010000001011011110110111110110000001010001000101111111100001011101010100010; 
out1756 = 128'b11110011000110010100101000110010110010100000100001000100011001001010001100100101000001111000011001000111111101001011101011100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1756[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1756, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000100111010010101101101010010110111100110100001010000100111001101010000011100100011101011011010011000110101111100111010011; 
out1757 = 128'b01010101111110111100011001011001000101000000110101011110110000110101100000011111000110010010011011011010111000011100010111111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1757[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1757, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110010011001111010011001110101010000011011000100101111010001010010110100010011010100101001101100001001111110110100010000101; 
out1758 = 128'b01011111001001101000000001111010010101001000101101101000110001101001011110000010110001101000101111100100110111101011101001101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1758[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1758, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110010011110000110010010010010110000011000001100011101010111111001011101011110110010001101101111110001110011110001111100010; 
out1759 = 128'b11011001101100000100010000100110111001100111010110110110010110011101100100100110111111110101100100000101010000100110010000101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1759[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1759, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110011100001011000111010100000110000001100000001111001010001101010100010110111010101010101110000100011011001100100011011010; 
out1760 = 128'b11010100111100111101101110000011000111001110111100001111000011101000101110111111101001111000100101000110110001001010101110111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1760[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1760, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001111010000010100100010111000011001101010110110100111110001101111010101100111000100100000110101110000000001110111001101001; 
out1761 = 128'b01101000001011111111001100110011111001101111110010001110010001110011001101011110111110100001000010111100010001111011101000101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1761[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1761, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001110111100000111101101111101110110000011101100101011110110100111101000010101011010011111000001111110110011001111101010111; 
out1762 = 128'b00010100100101100011011111111011111111111000100010001101001111111110010001011001011001000010001001110110111010000010011110010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1762[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1762, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100011000011111010101100100011100000000000010101110011110000111110100101001001100000100110111101010100011110000010011100011; 
out1763 = 128'b10000111001101111111110001101101000101010101101100001001011011000110111000101000010111101000011111110001000010001111000101011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1763[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1763, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001010010011011100110000100011100100101010000111100110101101100101010000100010010110001001100010011111000101000011010110000; 
out1764 = 128'b00010001111010010010011000101101011111101101110001001110110001110011010000010001010110100101011010101110101011001000000111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1764[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1764, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100011111001110001110001100011011111111111011100111000011011111101001100110010000100111101110101100110101001100011010010100000; 
out1765 = 128'b10110000000001001001101101101111110011000010010001010110011001101101100001111001111000101010110100000011000000101101000110011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1765[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1765, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110101011100110001000100011111010101000100100101001100110110010101111010011011100000011000101011000000101010100110000010010; 
out1766 = 128'b10110010010010111001000111001110110010011010101101001001110011100100000001010000011000000111110000101001010100101111111001110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1766[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1766, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111010100100010100101000101100001100110111101100010000101010100010110111101110000111010001110010100101011011101001111011001; 
out1767 = 128'b00111000000001110010101001011000010100111000110101110010110100101100101111110001001100011001101101001011110110000011111000101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1767[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1767, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010010001110101111110001011111010101011011110011100110001111101101000100010101010001111011110100011110000010001000111101111110; 
out1768 = 128'b11110011111011001110101010100101010011001111100010011110010011111010010110010100001110110110101010100101101101011011000011100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1768[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1768, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000101011101101110010001110101101111101001110000001000100011011001001111111011011000000010111111100101100010101110000011000; 
out1769 = 128'b01011010111110110100111111010001011001100010100111000101011001101110000110101001101011000010100111001110001010101101001000110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1769[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1769, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110101110010010101011110110100100101010011101010110100001101100010001101110110001111110100111001111111110111110101100000101; 
out1770 = 128'b10111001010010110111010001101111110010110011011001111011111111000110000000101100010001111000101001111010101111011001110100011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1770[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1770, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000001111011111110111000010100100101010000011001010010001111011100100011011010000110101010100110010110010001010100010000101; 
out1771 = 128'b11100100111101111111001101111111001111101100001010111011000011010010100010100000111110101110101000101110000101001111001010010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1771[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1771, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011100101111001111110010110111011001100100000000101100111100000011101000111111010000011000100101111011101001110100010100111; 
out1772 = 128'b00111101100100101100010000000010011111110111111010110001101010110000011110110001000110000101111100100110011001101101111100010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1772[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1772, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101101111010000000101011011011101010011001011111001001110110011011001100111000001101110001011100000100001100000001101011111; 
out1773 = 128'b00111111010100010111010010110110111101000011100111110100111110010011110010100111010101101000001001100000001110010101100110010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1773[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1773, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110000000000111001101010011111001111101101010010111011111000100011110011011110011000111000011110101111010001110111000001111; 
out1774 = 128'b10111010110000010100100110101001011001100001000011100001000101111001100000001001101111001010111100010000101011111011100010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1774[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1774, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110100100010101000111101101011100011111110001010110101010100011110110001011001000111000001100100000111011111011000111110001; 
out1775 = 128'b11011011011010000100000010110111011010110101111000100011011100101100000111011111000010111110010110110111000111011100000010110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1775[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1775, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100101010010011111100111101110011111101110111100100110110010001000010110110010110111000011000111010100000110101100011010001; 
out1776 = 128'b01001100110101011100011101110100011100000101010101101000100111010111100000000101000011101001011001110101011100001001010101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1776[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1776, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111011101000100101011000111000110000111111100001001011011011011110011110000000011010110111110101110010110011000111001111001; 
out1777 = 128'b11111101011001100101111110111010001111100100111001100101110010011101100010010110001000010110000000101101111001011110110101011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1777[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1777, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101010011010111100111101101000000010101010100010100110001001100100001110001001010101100000000011010100100000110001100011110; 
out1778 = 128'b11000110101111100110011000001001111000011110111110000110101010000011000100001101110110100111011100011010100011011111011010001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1778[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1778, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001010110110011111001101001110011010111010011001000111111011000111100010101101001011101110000111100100100101110001011101001; 
out1779 = 128'b11001001100011001100101000101111001110110110000011100001100010110010001111100100011011101001101010111111011101011111010000111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1779[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1779, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100000101101000101111111111110010101111011110100100100001100110101110010010100111010000101101001001101111011100001011111100; 
out1780 = 128'b10110110001010100010111100000011101100100011010001010101011100011111000001110101110101011011100101000000001010111011101010010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1780[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1780, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011011001100010000111001001010010110010001011111110110010101100100110000001001000011010001111101101101011101110100010000100; 
out1781 = 128'b01111010010011111100011110101000101001010001001111111110011101011100101001011001010110100100110110101111111011010011110000010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1781[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1781, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001101011010101101111000111100000001101001110011111011001101010100111100110000101110011001100110010110100010001011000010011; 
out1782 = 128'b11111000011001100000101111101001011011110111110010011100110101100000100000111111101000011110110111110001010110011011011111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1782[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1782, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001101101110000101011101100110100001010010001010110111110000011110011111110111111000101111011001111001011000100011100001101; 
out1783 = 128'b11111111000110001010001001000110010101001110011100011011001011010000110100001101011111111000001100100101110000001011001100111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1783[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1783, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000100101000010011111110011000000101100000011100100110000001100000010101100010001111110010011111011100111000101000011000011; 
out1784 = 128'b00111001001001101101111000100100011100001100110010101000001100100000010100010011110010000000100110001100010011110010011101110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1784[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1784, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110101010010100110101001111001011000101010000010111000101010001101001110111101101010000100000000111110011001011101111110111; 
out1785 = 128'b10101000100011111011010001010001000010110011000110001000011001111111111111001111000011111101100111001000000001111100111101101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1785[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1785, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001010110111100010011111110111011111010110011111011011001100011011101110101011000100110100000001100101011001111000001110000; 
out1786 = 128'b00111110100010110001111011111111110010000100000001000011111000101100100100001011111011001011111101000001011010001010000100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1786[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1786, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101001100110101001111111111000110101111111001001111001000011110101111011111000001001010100011000001110110011010000011011100; 
out1787 = 128'b10100101001001011001010100010000110111001010011100110110001110001111111010100101010010111101101111001111100011110111111001000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1787[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1787, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101110101100111010000000101011111000101010111101000111101110100100100000110011111110101100011100011100000001100001011011000; 
out1788 = 128'b00110100100101011111011110011000110011100010111101001010100101110001011111110000010011100011110001101000101011100110100100100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1788[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1788, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011010101111000100101110000010101010010000101001010100001010011100100101111011011011010101111010010111110010001100110111101; 
out1789 = 128'b01010110001000000001111110101110011101100010000010001000111100111110010111001111111100000110001101110100010111101101010000101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1789[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1789, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110101100001001010101101111001111111011100111101011100101000000110101101010110110011010011011011100100010110111000100000010; 
out1790 = 128'b01011100010101011110100010101100100000010010000001101010101011000101101100110011000100110011011010110000111001101111010111111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1790[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1790, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110100010001111010001010101100001101101110101111100101001000000000111000011010001101001101000001110010010001111011010010001; 
out1791 = 128'b10100111110010111000100010001011110011111101001011110101110011111010010000101100110110011011000100101110111100011111101000011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1791[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1791, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001010101101110000001010100110010110110111010100101011101110111010010000101101110001100000000110101111000000110101010111110; 
out1792 = 128'b01110001011011010011111110000111100111001000110111111000010110011111001110110011111011000111110111000000010101011111001100000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1792[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1792, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110000000001100010111010010110100010001011001010110001000111101000001011100101010000011010111100101001001000000101111010111; 
out1793 = 128'b01011111010110011100111001000001000110001110110011101101101001111000101011000010110110010000111000010100111101001010011101011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1793[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1793, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111100101111100000011011110001100111101100000110001101111000001010100110000111100100000110111010110101011011100111010111110; 
out1794 = 128'b11111100000000100110000000010011010111111110111111100100100100000001110111011110001011100100101100111110011001101000010110100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1794[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1794, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111110011000100101011110000001110001110000011010011000111111011101001001111111000011001100100001001101101010110000111110110; 
out1795 = 128'b01011000100011101010101011001000101011001000011101001101101101001110011101000111000111100011110111000001000001101010011111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1795[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1795, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000110110111001010100111001111001011001001100010001000111010100011001001111100110111111001101110101110110101111110010001011; 
out1796 = 128'b11101011011111010111001000110100110000110000100011001010010111111011011101111011010100110010000110111110000011110000001110011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1796[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1796, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101011010110000000101010100110110111010110101111001100101110111100101110111011101111100100110010000011101001000101100100010; 
out1797 = 128'b00101001111001101111010011110001001011000000111111000101100011100110011001101100100000011110100000100011111000010010111110011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1797[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1797, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011011111000101010101000001001100111001001100111000101110110100110110111111001111000101010000001001001011001111101011010111; 
out1798 = 128'b00011001100100110000001111100101011010011000010011100010100100000101000101111000000011111010110111000110110101001111001111111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1798[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1798, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010100000110100100100100110001110010111110110110010010000010111100001110110101000111101000000101011100001100011100001000101; 
out1799 = 128'b01000001100100001001101110110100110111011001001011100000110101111011100101101101001010111000100101101010100010101001111010001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1799[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1799, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100101100100100100011000000000110101000111001011101010011011111110000010010001110010101100011010101110010110110011110101111; 
out1800 = 128'b11101010100011100011100010011001100011001100011110101001111110100110001110110101110101011110001010000000010110100011011111000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1800[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1800, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101010110110101011111011010110000111000011101000000110100101101011110111000001010110000100100101111001011101010101010011110; 
out1801 = 128'b10010001001110100100100000010000000110011100001011110110001011000100011110101110010101000100100000100011101010000000110101001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1801[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1801, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011101010011011011010110111100101010011000111010011111010101010010001001111101010001001011001100101000101000101011011110100; 
out1802 = 128'b00011100010111001101110111010101101110100010001011011000011001011101100110100111011101100010110001100011101101000010011110101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1802[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1802, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110110001100110001100010000111000111011010011110010100100010010000110011100000000000010011000101111001011000001100111101101; 
out1803 = 128'b01001110101000010000000111001110001011011111100011011110101111000001111110001101100100111111011111010010100001110110100001001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1803[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1803, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111010100001001010101001001110111111000011111101011111101001110111111000111111011111111100110001010110011110101001000010111; 
out1804 = 128'b00000010110111101000010100011010101111110010000100110111111011000100111001110101100000011001101100101000001111100111010101101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1804[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1804, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010010100000001111001111000101000011111001000100101000000101010100011100110011110000010001101001011001011011100011001001111; 
out1805 = 128'b00100100101001000100011010110110101000010100011110100001100011110111011110011011111111000001010000001110000110000001110011110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1805[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1805, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001001000000000110110000010001011011000101010100110100011010100000111100111011101110000000000111010011001001111000101101000; 
out1806 = 128'b11001111001101011001110100000001100001100100100001100001000000010011011010110100010001100010100100001010001100100000110001101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1806[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1806, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010000111110000010010001110110000100000001001010000101011110011101010110110111101100101001101000111011100001001101111101101; 
out1807 = 128'b00111000000010001010000110011110110100110000101101010000000100110100110011011010110111001000101000100111011001111000101011110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1807[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1807, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010111000100110011011011001100001101100110000100010101111100010001001001010100101101110101101101110001110000101000101011110; 
out1808 = 128'b11110001001001001101101111001111011010001011000100011101010100000101110111000010011001100101101100101101001000111011110001110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1808[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1808, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001111011111111111001000100101000011011110000001111010110101001000110100000111111101010110100001101001110111011100100110000; 
out1809 = 128'b11101011000001001101110011111001011010010110001100010100000010010111011100000101110000100011001111001010011110010011001010011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1809[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1809, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001010110011111011000001100110000111000111101110111111010111101101101001011100100001110101101011111100010010110101100110001; 
out1810 = 128'b01111110111110100000101110001101001100110100110011100001110100110100101100011011010001000111000111111111001010101010001100110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1810[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1810, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000100101101100110110100110100001000101101011010111100100100001010100100101000000100101001100100111100100010000110001100001; 
out1811 = 128'b01111110011110010110101111001010001101101000110111111011011101000110110001010011100100100010011110110101010001110110011011101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1811[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1811, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110110011001101001111110011010101100001111011011011010000101111110100010111010000011111001001011001101011100001000100011100; 
out1812 = 128'b01100011001000001111100011001101100110010000111011100111100001101110111100010010101100100100001101011111101011011000000011100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1812[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1812, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001000100100110110001011010100111101100101001100111010101101000000011010010101100000010001001110100000101100110000100110000100; 
out1813 = 128'b10101000010111010001110110000010011101110010011011010001011001010101111110100011010010100100011010011111010010101001111000111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1813[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1813, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100010101001001110111111000100000110100000001000010011100100001101101111101010101000000110110011100000011010011001111110100000; 
out1814 = 128'b00000010101000000111000001001110001110110011111111001111001000001101111001000101000000010001011001001010010100010010100101010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1814[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1814, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000000101110100010010000011101011010100011000111010010010101011000111010111110001111011000111100111000100111011011010110000; 
out1815 = 128'b00010000101000010011110110001111001110100111111011100110100011100010100011111110101101000101100100001001100110111110010010010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1815[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1815, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101001110000001110111001100101110100001001100010010010110011010110011110111011110111110101111011011001000111010101010111101; 
out1816 = 128'b00101101010100000111000101010000011111001011000100111000100001111100111100110101010001010100100010001001001101011001101010111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1816[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1816, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011010110000010010000100100001100101110000100011011000001111011110011100101101001110111011111011011111011111010000010111000000; 
out1817 = 128'b11111100010011110101001101100000001011100001110101101110010101111101011100001110000101011000101000000101001111001101001100111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1817[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1817, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010101100011101011001111110010100011110110111011100100110001000100010110110100101000110001010010010111110110111110011101000; 
out1818 = 128'b11110101110000111110010100110101010101100010110001111111100101010011001010101000001110110010010000110001100110101111101001100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1818[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1818, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000010010011011100001010011010001001110001110000111101101101111110100010001100100110000100001101111111101000011101111000010011; 
out1819 = 128'b10001010011100010101110101011001110010010010001111000101111010110111010000000001011101111111100100101100111111001101111010100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1819[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1819, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101100101111001111110001111010000110101010110101100011010110010000001011011110011010001011111011000100110000111000111011101; 
out1820 = 128'b01000000011110001110011110110000100011011010110111010100010101001011111010111011000110001111010010100001101110101101010010111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1820[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1820, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010001100001010001011000000101011000000100000010011001111100100111001011111010001110110010001111100001001010001100101001110; 
out1821 = 128'b10110100011010101110111111101010110000010101010000101011101110000010011010111110111011110010000000010001100101010101110110001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1821[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1821, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101010110011100101100011010100110000001110100110010001010010111110100011101010100100100010011100001001101010110010101110001; 
out1822 = 128'b10010000101010101101000010101110101000000010111001010110111101101010101110100110101010111000011111100100010000000111010110110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1822[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1822, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110101111101010100000101001110110101011100010010000110101000111010010010110011111000101011101100111001010010001101111111111; 
out1823 = 128'b11001110001010100001011100101000011110011011010110101000101001001010000100100010001001011110010011100111101101111100010001110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1823[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1823, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001111100111100001100100101011111101100011011111000100101101111111101010101001001001111100101101000110100100110110101110010; 
out1824 = 128'b11110010101101010011010011100110000001100000101001001010001101000000010100000110100001000000000110111001011001100010011011110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1824[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1824, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011011101001111011001011000010101010110000010110100111010100111110011010101101111101110010001000111100111100001011100100011; 
out1825 = 128'b10000101010011111101010000000100010000100000001100011000001010010110000010100011010110011001100011011010000001010101100001111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1825[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1825, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000100001101101000110011100001100001111001011111000111001110010110100001010011000110000100001011101010110100100010101000101; 
out1826 = 128'b11011001010010011000011100111011010100000010111000001000000010101010010111100000110000001000100011001010111111000011100010100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1826[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1826, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000111111100010010111001110111011000111101001011100111100000110010010101011110001111100110010101000100111111010010101000111000; 
out1827 = 128'b11101010010110110100000100111111000101110011110011110011001000100010010011111011001110111111100111101111011100100001011010101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1827[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1827, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000111101100010100010100111010110010110001001001101111000110110111001011110111100110000110011101110111000010101101010110010; 
out1828 = 128'b11010000111100111110110000100000000011001001110100000100111001111011000011101010111100100011000011110010011100111100001100111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1828[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1828, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011011100010101011100110110101011101111000110111010001000100111011110000010010011000010101001100111011001010001110111111110; 
out1829 = 128'b10011100010010100000011001110001000001010010110110100110111001000111111101011101001111000010111110010111110100000000011010000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1829[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1829, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010010111000111100001100000110000110110101010001110000111000100101011001011101010010000110101001101111010110101111101001100110; 
out1830 = 128'b11000010100110011010010000101101011000010010100010000011111111100000111111001010100101111010011010101001110111011001100101111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1830[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1830, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010101100110110100101000110101100101011000011010111010000100010010001110100000010001011010110101011010011111011111110111111; 
out1831 = 128'b00100010011100000111111000111001101010010001000101010101011001110111111001000001101100101010111000111001111010101011010000110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1831[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1831, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000001000110100101011101010011011001111011010100100110100101010101000000010000111111101000111110001101001000101110111110100; 
out1832 = 128'b11110001011111111101100101010101111111101101001011111001001101011010011000011010101100000011101001000001000110001010000100100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1832[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1832, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111110111000111000100101100001010111100000011110011101100110100001110001000011010101100001100111010100111110100010100101000110; 
out1833 = 128'b11101101100100110000101011100111110001100001010100011010011100111011010101111110010011100011100100010100000000001001111011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1833[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1833, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100110100100000000101101011110101011001111110111110110010011000001011011101101111010010100111010110110010101101001100011111; 
out1834 = 128'b11011111010100000100010101110100101001101110110110000100000100000101000110100101101110000100001011100000010110010011111100001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1834[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1834, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001101010011001011101000110000111111100100001000111110100110101001001001101011010011011111010100011010111010110000111101011; 
out1835 = 128'b10101001001101101000101111011011000000101111111000011110001110001001101101101111010111100101111100111100101101000010110100010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1835[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1835, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001110010100010100101001100010010000001101010010010001000000100101100000101001000101011101101100101011001110001100001001000; 
out1836 = 128'b11111010000000110001001000101011111111101000100101110011111001110000010101100011000001001101111000110011110001001101100101011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1836[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1836, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011011100101010001110010000101011100011001001000111000001100001001000001101110110100010100011110101110000110000111010000111; 
out1837 = 128'b10000011100001000111110000011011101010111001010111101100111010110100000001010100111110011111101100111001100110001110100111110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1837[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1837, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111000110001010010011111111101101000101000100110101101010101111010011101101101111111011010000011100111110111100110100101001; 
out1838 = 128'b01000001011111101100000001000110000111111001101011000110110010110100110001000101100010001011001101111000111010100010101000110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1838[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1838, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010111110110101100000000111101100010011001110011100111101111011110011001101000110101111100001000111100001011101011010100111; 
out1839 = 128'b01001100011100101010000100010100001101110001100001001100010000000101110010101101111111101111011110111110000011000001111001101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1839[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1839, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111001110000100110110100000001111011010000001110011000110110000100011101101111101100000101001001001101101001011111110011101; 
out1840 = 128'b11100011010000101111101000010110101111111100001010000101010110111110110110001101100010000000000010000000110101000110101010000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1840[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1840, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000101010100110100001001001111110100000000110001101001010100011110010101011011110111100000010111011011011110111010101010011; 
out1841 = 128'b10011010111111011101000111011110111001110011110111111110110010011010001000000101011000011000011111000010101001011110000011100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1841[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1841, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111110111011110001000100110101010001001001000100000001101010111001000001100110000110000001010100101001011100011100111000001; 
out1842 = 128'b11111100010110001101100001110110000001101111100101010000101100110010011110011001110000001111000110110111110010010010100010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1842[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1842, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110010111111011000010110000110101111100000100011001000110101011000001011010010011100011110110001001000110000101001011000100; 
out1843 = 128'b10100001110111010100101001010001001011101110110111111111011110101011100101100010110011000010000110000110111110111011000111110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1843[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1843, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101010010101100111101101010011110101110000100101111011001010110010111101110010000000000110101111101101011011001001010111010; 
out1844 = 128'b00111110111010011010000110111110010001001110010000000110010011111001010111000011011010010010111011101000011001011101100011001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1844[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1844, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111000011101000110110100100011100001110101000001010101100000011000000000100111100101010111111111101100101110111101000011111; 
out1845 = 128'b11001010000011010001001101011000100010011110110001001010110010001011101111011110101000100101101001101010000010100010101001110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1845[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1845, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011101011110100010000010111110011011110110101101101110100010111111111110101010010001000001101100100101101100011111011101000; 
out1846 = 128'b01100110010011000100001101110111011011111111011110111010110001100111011110111111000111011000100111001100011111110110110101010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1846[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1846, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101011000101101101100111000100110011001110001010010000011000101001111110000100110100110010100010100010111011010100000000000; 
out1847 = 128'b01100010001010100111101111001011010010001101111100001010101100011100000010111100111100100100110011100001000011010001100111111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1847[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1847, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111100011001000111100000010000000101010011000100001001000011100100000000110110100110011101110100110010010110001110001010000; 
out1848 = 128'b01111111000101100001001001001101010011110001011101101000111110110001110101001111100001110001000001000111101110101110100000001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1848[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1848, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110000111011100001000111110000100011010000010001101100001100110011001001010111111110110101101111011010010111110000101011001; 
out1849 = 128'b01001101110001010010001110111110110111100000110000111110100000101101101110000101100011000001100010101010010111100011101010110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1849[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1849, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000111111101011010100001110001010011110100100111011101100111111100011011010010111011001001001100100100001001001101111111100101; 
out1850 = 128'b11100100000111100000010001000100110001000111000100110000101101110111100101001011100110000100101000010110000001001010000100110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1850[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1850, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101000010100101110111001110111111000111000010011111111000100000001000000110101101101010101011000011000010100011111111111000; 
out1851 = 128'b00101100101111100000010100110000001100100111101001001100010011110001110111000010000100000000000111011010110011010110001010100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1851[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1851, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011110001001110010001010001000110010010000011110100010100011001011000111110011110101011100010110000000111001111010100000011; 
out1852 = 128'b10110100000001001110000011100111001001110100100100101111010000011010111110001101010001111100000100110100100011010110000000110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1852[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1852, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001111111100101111000001001010011000001001001110010010011010110110000011100001011000100001110010010000001000010011100110010; 
out1853 = 128'b11001110101110010000011101000111101011001110110000000101011101010100010001110110100000000001001111110000100011110010000110011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1853[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1853, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101000101010110110000111110110011001111101111000010000011100010110101010100110011111010100000111110110101111010011110101111; 
out1854 = 128'b00001101010000110010100010100110111011110101100100001001100110000100111111110110010101110110001101010100111110011111110011101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1854[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1854, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001011110000010011111110100101110011100010101000100110110000010000110001100000001011111001000000010010100111100110010001000; 
out1855 = 128'b10110001001010111110010101110011010011010000011110100111101111111000111011110101010010001111011100011011001010001011111001110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1855[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1855, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011101110111110010011110000111011000100010001101110010011110110001000110110111001101100001000001110010001000010100010010110; 
out1856 = 128'b11101000011110101011101011111111100001101000101000111001110101110101000101011010100101100000110010111101100010011100001000011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1856[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1856, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011100110010010010110100101111110111001110001011100100100000010101101001010000000011111110100101101111000010010010100000111; 
out1857 = 128'b01011110110101110001111000101111101000000100001100110011010101000100101110010011011110100100101010100001101101100101001010101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1857[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1857, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101110010001000010111101101110111010001101111011100001111100110011010101010111000100000000111011001011110000100110011100101; 
out1858 = 128'b11101001101010000010000110010100101010101111110011010110100100100111000001101000011101001010000000011010010110011001000111010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1858[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1858, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010111001011111000000100110000110001101001110101010100111110001111010111011110010000111100111101110100010110110001110101001; 
out1859 = 128'b11001111000000010011000001101001011100101001100111011101001000011001001010100100011100110010111011101111101110001111001001110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1859[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1859, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011010010001111011010100101100101001010111110010010100001100001001010010101100010011100110100100000100111111111101101100111110; 
out1860 = 128'b00111100001101000001010111101001101010000101100100101000100000010110000111101110011010110111000101010010100110000101001000111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1860[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1860, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101000011001110101100001000010010000000000100000010010000011111011110101010000101110111101001000001001010101010110101010000; 
out1861 = 128'b10000110010110010101001110111111111110101000001111011110100001110000000100001100110101010101011001011100100110111011111011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1861[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1861, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010110011010010010101110010101000010111111000000011000110000001011010011011101010010110110001100100010000101100101000010100110; 
out1862 = 128'b01011000010010111100110000000001111001000100110101101000010110001010010011101110100101111110110000010000011001001011001101011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1862[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1862, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101100011101011100010010010100011011011110000000011011001010001101111110010110101100111100001111001110000001011110000101000; 
out1863 = 128'b10010100101111101110001011111001100000010100000110111011011101110110100001110011101110010100000100111001111001111011101101000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1863[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1863, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000010100001001011001100000100100110100110101111111000101010000011011001010000011001001100100111011011010010101111100011101; 
out1864 = 128'b01000001000000111111100111101010100100110000000100000010001010001000100010111110000011001100100011001110100010100101001110011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1864[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1864, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100001011001101010010010001100100110100000100011011110101001000001010110001100000001010000111000010000100010010010010111100; 
out1865 = 128'b11100010001100010010000011011001010101111001010100111100001110101000001010111001011111000001001000110110000101101001011101010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1865[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1865, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110101011010000010001000101100010001100001111010000110100001010111111010101011010101111011111101111111111111001000111010110; 
out1866 = 128'b00000011001001000100011001110100111010001011110011110101110101011100011011010001100001000110011110001101011110111001110011111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1866[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1866, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110110110011011110111001011101110010011000000000110100110110100110011111100010110110001010110101010100110100010110010111010; 
out1867 = 128'b01110100111111110000001010110110101011011001011000100001001100011111010011100010100010100010110011011110101111111110010011011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1867[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1867, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010000110010001101011101000100001011101100100100110011000101100011110100100011101100011101011111111111110011101111010100010; 
out1868 = 128'b11110111011011110100000100001010111000101111001110100110010100011011100000000011101011111111110010111111001110010001111000001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1868[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1868, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110101100111110101100000101010100110100101101000010010011011100101010101000001101000000010000101111000000100000111011110110; 
out1869 = 128'b00001100000101110001100011111001000110001111000011110000110011101011010110000101100101010000001110010000111000010010110101000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1869[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1869, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010110001000010010110001111011100010101101100011001000000100001111000010001110110110101010101100010111001110010100000100110; 
out1870 = 128'b00110111011010110100011110111100001010101011111110010100101010100111111000000001100101110100100101100011011001010101010100101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1870[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1870, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100000010101101110101111101110010110001000011000111001010001101110110011011000101100010001000011001000011010011110010010000; 
out1871 = 128'b00111111010100110001010110010011001111100001011101111001101110011100100101010010001001100011101001001001010111011101110110011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1871[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1871, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111100001101111011000001111100111001101101010010001100011010111001001110010110001111000011011111010010110000111000110000101; 
out1872 = 128'b01000101110000100100011011010101110011001011011100000010101010010101100101110101000001111011011101000101000101100001101111111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1872[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1872, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011001010001110101011110011110100001011101101011000001111110110100001011101101100110110101100000100010011001111111100001101; 
out1873 = 128'b11100011100011100101111010010010100111110010000011001110010111000110001111110110110010100101110000010011010010010111100100010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1873[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1873, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111001111101111010000010110111000110001110000010010011101110111111110001101010110010010011000100000101101010100010101100011010; 
out1874 = 128'b10000010011111100010110111011000011110100011100101110010111110110111010110100011110010111000011110101011011000111100111000110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1874[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1874, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001001001110110111000110011111010011010011111100010000011100101110010101101100100110010011101010111010101011000011010101010; 
out1875 = 128'b00100011011010111000010111001101001100010001001100001111001100001000011101100110111110101100010110100010101010001000010110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1875[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1875, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001101001010111011011101101110010100001100001010000000010001100110110110000010011000010001100101001011100101010100011101101; 
out1876 = 128'b00011101100000001011001111011000000001111011101101100110111010101110011001101110010101101000101010111010010110101001000111000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1876[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1876, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011100011001010111100000001101010111000001010010010100000001110110010001100001101000101000000101011111010010000011010101111; 
out1877 = 128'b10100100101000111100110111011101111100001101110010011111101110011000011001010111011110010111001010011111110110011001000100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1877[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1877, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101010010000110110000000010101010001111101110100010011011110010011010010001001000100100101111010110010010100100111100010100001; 
out1878 = 128'b00100111111011111100001100110100100110100000000111011010111111000001000101110110000111111110110100100100000110100101011110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1878[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1878, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000111110000111101011100000111110110100110011010111000010000011000110110011000111000000000000111011100110100001100010001010; 
out1879 = 128'b10001101000110100010000000010011001111001111110111101001100010110000110110101011010001101101010001110100001100110000100100101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1879[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1879, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110100001100100101000010111111100000100101100101100101010111011111011111110011101001000100011100010011111001001101110010100; 
out1880 = 128'b10011001010101111101101010010100001111101010011010001011010110101111100101110101000000100011011110010111001101001101001101111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1880[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1880, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011100100111111010001100100100110001000111010111101001010100001111101001000011001010111001110001011000011011011011100001101011; 
out1881 = 128'b00010001111111111111100110110011010000001011011000010001011100110010001011001100110001111111000100110101110010100011001110101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1881[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1881, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100011101010100010100011010011101011101001101111011100011011101000000000010000100010001000001011101010000101011101010110110; 
out1882 = 128'b01110001100000111101001110011101110111010110111000011001000111110111000011010011100110111010101001010100011000001001000100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1882[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1882, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011000100101110010100101110001010110010110001001010101001010010000001010100010111100011100101110001101111111100000111110110; 
out1883 = 128'b10010110011001011111110100010001010111111101100110100101011100101110000110011000000111111100100001100001001000101101111010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1883[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1883, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110111011110101111010111100000001100000010011000111100001111001111010110010010001100111001001100101110001000111000001000010; 
out1884 = 128'b00100011001101011000101011101100010110110100000000011000110101010000000100000100010010011001111111000011010010010010110010111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1884[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1884, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111011010101111001110111100110010010000011101110011000110101000000111100110110110011110010011111100110100101101001001101001; 
out1885 = 128'b11110101101001011010010000111110100100111101111101010101101011001111000111010001001111000111110111111001001000111111001010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1885[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1885, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000110101100001101101110011000111010000010010110000111100110011111001111110101010101001000100110011111010111011000110010010; 
out1886 = 128'b01100110101100001111110110010110010110001111110100001110000000110000111101011110110011011011101100010111011100100101001000110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1886[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1886, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110010110011100010010110111011011110010101100100011111011111001011001001100000000000000100010011100001100011000010011111100; 
out1887 = 128'b01000010001100101011111011110111011100001111111111000011010001001101100001001110001100101110011011101101000010011011001100110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1887[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1887, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111010010010100000111111110011000101001010110100011110110000110111000110010000001000011101000011001010010011111100010001001; 
out1888 = 128'b10011111110101100101101000101011001101110000100110111111011100011100111011010101100011100001101100010011111101011110101111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1888[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1888, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001011110101110110110010011000110010101011011001110011111111011010110100011010101000011000101010111010110111100101011010111100; 
out1889 = 128'b00001000101100000011100000010100111001011111011010011011110011000111100110110100110000111000001010000000100011100110100111100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1889[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1889, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000110011100110110100100110010001100101111111001100011100001011111000001110111110100111111100101110010101101100000100111101; 
out1890 = 128'b11111011100011100011111001010001010010100100011001000010011100100111001110101110110010100101010010101111101010110101111111011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1890[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1890, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100010101011000110000011011010001101001101110010011000000010110111110110111011010111100001011110111010000101101100110011101; 
out1891 = 128'b01001000001110101001011101001011111001110111000100011101011010000010001110111011001010001000011110011010010100100110110110000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1891[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1891, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100011101011000100100011010010111101111010101010101111001110100111011010010101011110000100010111001011100001101010010110000; 
out1892 = 128'b11000011000000010110001001010111101111011110000110110110010010111010001100101010001010110001100000000101110110110101001110111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1892[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1892, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110010110010101100100111100100100011111111000000100001100011101110101000000001111100000001010111001110101001100110011100110; 
out1893 = 128'b11000000101100011101000010100110000000100110001101010101011110011011011011110100000111001111101100100111001101000111001001111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1893[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1893, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010110010011110001001110001100100000101000011111100001001011100110110000101111011111101011010001001001101111001101100010101; 
out1894 = 128'b10101000111111110011101110100000001101101110011110010111001111011000110001101100110100101111011101110100110101111010010010011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1894[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1894, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010110101111001100010000110110000000100010100000001011001010111111011001110110000001110101111001010111101100100011101001011; 
out1895 = 128'b00101001000110000110000110110110000111010000100011100101100100100110010100111100001010111011111001111001000000111111000110011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1895[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1895, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000010011010111110010010101101011010110100110010001000100101110001110001001111101111111011010010011010001001111000011100100010; 
out1896 = 128'b01101010000000110000111000101100111000111100001011010011111010001111001010011011111000100110100111110001101001011010111111111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1896[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1896, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100111100101011101111000100010100101001110110001111011011011000001101001000010001000100110110000101110110011111101101111011; 
out1897 = 128'b11010110001000100110000110111010110111101000101100011001001000110010011010001110001001100101001101010011100100000111011011100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1897[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1897, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101010111001111100101010110100000001100101011001101101011010001110101110111111000101010111110110111101001011011111110001111; 
out1898 = 128'b01111101001011101111111110110011111100011100111011001000110000111110010001111001000110100000001111111000010110110011101100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1898[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1898, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101100110011010101001010010101010100011000100101010010001110000110110111010100010100000100000000001110100011001110100010000; 
out1899 = 128'b10010101111001011000100010111110001011101000000100001000000011011101000011001001001111111001001111010010011101010011100000101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1899[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1899, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100011011110100100011000011011111010001011100110001011011111100111101111000101010010001110101000100000010000011001010110111; 
out1900 = 128'b10000101001111011100000001011101000000101101000011110011100100101111010101100010111111010000101111100010001000010011101110100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1900[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1900, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111110111111111010111101000110011111010001001101101100110101000110000000000001101101000100010111100011110011001100000010011; 
out1901 = 128'b00010011100011000011100111111110110010011101000110001011110110100011111001011001101000001001111001100101100000111010110010101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1901[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1901, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010011100110110101100011011101111010110001111101001110011000011101010001111111100110110111000111011010100100011011100010100; 
out1902 = 128'b11011011101100110111100111001001101000001000001100111110100001010100110001101011010110100011001100000101110000100001011111011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1902[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1902, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010010110001001010001111110011101111001110000101101100110010100010110100011010000011110011000001110000001010000011100001100111; 
out1903 = 128'b10100111000011000111010101010111010010100101111000001100000110001110010101001001001100011010111100011101101111011000000111111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1903[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1903, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101111010100110111100010101011110110011110011010011001101100101100001100111100011100100001110000001100110010001000110101000; 
out1904 = 128'b01000100111001110000001111101001000100011111111110001101001100010110000101010011110000000110101100101011010001111010111101011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1904[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1904, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001101101100000101101110111010101010101010110000110010000111001000010000100011000110011000101000001011100111110111011110111; 
out1905 = 128'b00011000010101111011111100011101110011101010001000100000011100110001100000001111000110010100100111110101000101110111101001101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1905[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1905, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001101111111110011101000010011111010001011111100100000000010000111111010101111010000101011100001100000101001100000101010000; 
out1906 = 128'b10000100100101101100001101110101001100011110101111100101000011110110001010000010011110011010101010010101001111100111000011011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1906[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1906, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011001101101000100101111000001110110111011100111111110100011110111010010101011100100010011110010010011111011110000001011010; 
out1907 = 128'b00010111010101110011010011010011110101001111110001110011000111111001111110100010101111100101110110011100110100110001101111011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1907[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1907, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100011001100000100010111011101010110110101111110011010000101010001100000001001000111101100111011010111000000111001101011000; 
out1908 = 128'b00100111100011101001001010010110111110001001010010001001001100001101101001101101100001111011110010101111111010001110000000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1908[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1908, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000101001101101101001000100000000000111010100001111000101110010011011101100111101111001001101101101001101101000010111111101110; 
out1909 = 128'b10010110001001011100011001000110110110111011111111110110010000010100111000110011111100011111011100110100101110101001000000000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1909[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1909, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000110010011000000111101001111000010100101111011101000010011001101000000011011101000010101010000101100001000000000000011000; 
out1910 = 128'b00101011001100100110011001001011011001011000011011001000000001100100111000000101110101010000000101000001101101100110110010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1910[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1910, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101010010010001100101010100100101100000010000101100101110000000100111110000010000101100010100111100011000011011111110010110; 
out1911 = 128'b11000001110001101000001000000000010111111111000011000010011000100111000100011000111101011011010110110000101111100100110011010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1911[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1911, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110111000100101010101111101001010011100100011010010000011110101011111110011011010010010101111101101110111111001001111000001; 
out1912 = 128'b01111111110110001000111010110111101000011010001000000000111101000010111000010011101011100001110000100010111001111100010100010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1912[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1912, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100000110101111011011001101111000100100011111000000011000111101010101000000010110000100100011011011010010110100110001101001; 
out1913 = 128'b00000000000101010001111001010000101111001010010101011110100000101110110111010111011100010111001010110001111101001000110101110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1913[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1913, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000100000111001110010110001000100011011001100000110101101110000010010111101100010000001000011000101010001010110111100100110; 
out1914 = 128'b10110010100101001100011011101110101101011101001010101111010100000000000011100110110011100010110000100110111010001011001011110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1914[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1914, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100100001001101000101010101110110010101001010000001111001100010101110000000100111011000010011011101110100110000110100100110; 
out1915 = 128'b10101000100110101001110000110111100011000111010101011011101011111100000010001111101000001100001011010001011011011010100110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1915[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1915, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101000001100100111101110110000100001001001010000010111110010010110110111111001000110011000101000111001001100101011010010101; 
out1916 = 128'b01111111011100000010101010001001101111110101101110010100101011100111000011110100110010110101010010011100001001111110101100011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1916[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1916, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011001111110101010110011110011011100011010110100011000010110000101100111101000111011000010011110001001111101111010111000110; 
out1917 = 128'b11110101000100100101001101010000011010111001101111111111100011010000001100000001001010011000010110100001101100110110101101111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1917[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1917, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110100001110101011001001110111110111000011010000011001110110010100011010111100101000000011000101000010100110011110010011000; 
out1918 = 128'b00011010100010001111110010010100101100110101010010000010101100000000111000111011001000111110001100011111001001110100010110011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1918[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1918, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110100010111100011001100011100101101001111001000001010111100110011010101100011100001000010111100101010010100110110100011111; 
out1919 = 128'b00001111101001011101010010111010101011010101001001010000001100101011100000110000100110000010101011001111011111100010010011001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1919[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1919, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111101100111101010001010111010100100111110111010010001011010100101011101010110111000100010000100100111110001101100000001110; 
out1920 = 128'b11111110101001100111110001001101000001010110101000101110101000110011110101101000100011000001011101011001110011100010100101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1920[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1920, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001001010010101001101110001011010101110001100110110111001001001111101010101100101000010000101111110110000110111100110111000; 
out1921 = 128'b01111100010001101001001101000001011100010001011111101000101111111010111011011110111111011111001000100000010011111110111010000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1921[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1921, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100101010010001110010001010100101000100100100010100011110110111001110100110000101011010000111001111111001011100101100001111; 
out1922 = 128'b00100100011101000111011000000101111100101111001011011110100011010010001011101101100111010111101000001100011011101010001101011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1922[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1922, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000111000010100000011101001011001100111110010011101101011100001000111001101010110001111100010101001001111111000100010111010; 
out1923 = 128'b01110110001011100010111001011100000101110000000000100100010011000011001001110000111100000100001100110111111101001101110001100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1923[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1923, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000000010010010100001000011001100001110000011111010110000101110010000010111100101101111111110011010000100110010010000100010; 
out1924 = 128'b11101011101110100101000100000000111111000010101000000010010100101110011010101100010111100011011000111010101010100110111011000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1924[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1924, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101111000110100111011001101001011101000011010000111110101110011100110000000101101010000001100101001000101110110100000000101; 
out1925 = 128'b10100000011100010010110111010111010110101101100110011010001010101110111001010011010101001000001000000001111100011000000000110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1925[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1925, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001101110001001101110000011110000010011111011011100011101100010110000101011110000111100010000010001111010010010001100100101; 
out1926 = 128'b00110100010011110000101000111110110001001110000011110000011111011110110101010101110010001100001010101010100111000100101101111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1926[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1926, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110010110001010001101110111111011111101010110111100100010110111011011110100001111101100110011000111110001000100000101110100; 
out1927 = 128'b11111000100101110011101101101110010011001100001011111111111100110000000010000001010111110101111101000101000111110101000111001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1927[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1927, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101101001100101100110011111100001000111011010110001000101101110111101101100010100100001011010001111011100101011100110110000100; 
out1928 = 128'b11000011010010011010011011011110100100011000001011000101111000010101010010110101101001100011010100011000001110001000000100000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1928[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1928, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001111011101110011001110110000101111111110000001000111011010000111011111001111010010001100100000010100001110101111000010010; 
out1929 = 128'b01100000101010101100110011110010011001100101110000001000101001111010010100101001100110111101011010100000000011001010001111101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1929[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1929, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000111110011001110101110101110101100000011110001101111001101001011101110110000000100101011110101100100110100110001101111101; 
out1930 = 128'b10111100111010010011000111110001100110111000001101110000000110010001001111000111001110000001011000100111001000111111011000010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1930[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1930, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010111101001101101010101010011001110001100011010101100111100011001111011000000000100010010011100111010111000011011110010101; 
out1931 = 128'b10000110111100000000000111011111000000000011110101000000011011000011100010110011000001111010011000111001110000001010100100101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1931[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1931, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010011100101000110100001101100001010101100001101100000111101110110100100000111010001101011100001011111111010010001101010001; 
out1932 = 128'b10010001111011101001010111111101100000101000100010001010001100011001011000001101001110111001100101010011011010110001011010100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1932[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1932, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100011001101001100000100011111110100011111001000011000001101111101100110100010111111011110111001011000011001100001101010100; 
out1933 = 128'b10011100010001011101101101010100100001101001101100011100010000110000000011101000011011011111001011001101000101000001011011011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1933[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1933, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010010011101100110011101000110010100111001100010011010000001111010110010011011001001100100010111110011010010000000100111111010; 
out1934 = 128'b10011111100010000111101101110000001000000011000111100011010101101010111100011110001011001001101011001000000101100010100101001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1934[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1934, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100011101000101101100111110001001010100111000111001110011011000101010000101000010110001000100100010100010100100110011011011; 
out1935 = 128'b11011010000001110101101011001111100100110110010110001111000011010010111111000011100001001101110111011101111011001100010001011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1935[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1935, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000000111101010001001011001000000001101110011000111000101010110100010001000011110111110010000010100010100000010001010000011; 
out1936 = 128'b10100000100110101100001110111001110010000111000110101010110100110011110101001001110000110001000111110001000001010001110111011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1936[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1936, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111100011101011011000010101101101000000001100100110000101101111011111100011000001001111000100100110011010100000001011001100; 
out1937 = 128'b10110000101010001101100010001110010101110110100010001000110001011010101110010010001111101111100000001001010111101101111000000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1937[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1937, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000110101000100101010110010101001011111110110000111011010110000110000101000100110110110010110000101001000011001000001100100; 
out1938 = 128'b10111001101011111101100001100111010011100011111001100110100011101101100001100100101011101011000101110001001011101111001111110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1938[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1938, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111010111001000001100001111100100100000000110010101010100001001101111000010100011010011010010010110111101101000010011101011; 
out1939 = 128'b10001111100110011111110101011100111000110100001101010100110010001111101011110100111001100101101000000011110010100110101101001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1939[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1939, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100111000010011000010110001001110100010101010101110011000110100011001010110000111110110111011111010001001000001110100000110; 
out1940 = 128'b11010110010111001000110001001101101010010101110011010010111110000000001101000001011101111110111011101110011100010101111001001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1940[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1940, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100110101110001100001011010011011101100000001100001001101001011111111010111000110110111101100101101011001001101110011100000; 
out1941 = 128'b00101010100100001101001010111000001100000001111001111110100110000101111000110000101100001101010000010100001111111101000011011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1941[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1941, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000100110000100101000000010100011101000001000111010001111101111011101100110000011110100101110010101101010011011111011100000; 
out1942 = 128'b00000101001000101111011011100100010110000001010010100010010000111111100011010110100100111001110101010101100010000011010101100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1942[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1942, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110011001000001111011001111001011100010010111101010011100001001011110000010100011011100110011111001000011010110110011111101; 
out1943 = 128'b11111111100010101011100010001110110011101010100010010110010000011000110000111110110000010110111000010110011100111110010011110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1943[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1943, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011011111110101101110011111111101011101011011001110101110111101110110010000011010001111100100110101111001101011011000010000; 
out1944 = 128'b11100010001111000111001011101000011100001010111101101001111000110011100010000000111010110100111100001010001100101100010001101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1944[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1944, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010110101100001110100000101011011000010110101011110000110100011100011111100100011001101001000100101101011010011001100101011; 
out1945 = 128'b00111111101001001010101001010011100111010010101010111001001001101101000001001010010111001011110100001011010011101100101100000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1945[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1945, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111001001101101100100001011110101111100100000110111110001101111100000100010101011101110010001111010010100000101110010001100; 
out1946 = 128'b01001010110111001110110110101110100011011000100100110010101111101011101000011111010101101001110110011110011101000001100001111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1946[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1946, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011100101100111101101101000011001101111011011011100010010011100011111110000011110101100000100001010110001010011110010001110; 
out1947 = 128'b01010100111100001110101101111110111111010111000101110110010110111011001011101110101100100000101010010000101111010110110101011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1947[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1947, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010011001000001111101011101001011111011000000011100111011011001101011000100010000100000001010101001100100011101001110110111; 
out1948 = 128'b10010010101101101000011010100000011101100000010100101011111100111000010000001100001001011100110101001101110011000011100001111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1948[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1948, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000111011010110101001000100111011010000100010001011111100011111100111010000010001011001110110010111110010110000001111100110; 
out1949 = 128'b10111100100010010100100011111001111101111001110011111000000010001100010101101110001000101001101011110111100110110111100010011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1949[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1949, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101011110111011000101111101101100100100011001100000101101001110111011100101100100010001100101100011010110101000100001101101; 
out1950 = 128'b01000001100101100011111011000010110010110011010100111101100111110010010001111111011110111101001000001100100101001101001100101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1950[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1950, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001010000101101110100000101110001100110100101100001000010001011111011001111110001001011010101110011001101111100001001100101011; 
out1951 = 128'b01001000111100010010100001001110110100111001010000010001011000111111001001000110110111100010100010101101101001001001100111011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1951[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1951, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101010011011001011101000100010001011001010001100011000100000100100011001000101101001000011010101101000110111101111001100000; 
out1952 = 128'b00101000001111100101100110111110011100100010110000011001110111011101101011100111000100111011011100000101110101010111001110110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1952[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1952, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010010100001001111000011000100111101100000110100101000000101010011011110101000000110011001111111100000001110100011001100111; 
out1953 = 128'b01101110011101000111010110101010011110110101011101000110100100010001101001100101010101100011000101100110111011010111010000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1953[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1953, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001110100010010011110011110111111101100110000010001100100000101100000111010010101101001000110111001100100111100011100010001; 
out1954 = 128'b10001000100011101011111110011001110110100100000001011000100011111001100110100000111000001101110010001100111101111010000111010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1954[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1954, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110110111111000110100101101110101011001001000000000101111010000011011101011101011110011011110010101101010000100011001011101; 
out1955 = 128'b01100110101100000000111100010111101101011101111001011110110001101001111000100101011000111110000110101101001100101011011000100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1955[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1955, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010000000011011111100000110000110011010001110011000000111010100100110101111000111001101100101110100101111100011111101000000; 
out1956 = 128'b01001011011111100101011110101001010110001010010000111000001001010010000010111111011001100001111000010011101111101101100001111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1956[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1956, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011011000000000101110100000111110100011110111110100001110001001011101001100010110100000001001111011010010101011010111110010; 
out1957 = 128'b01111111111110001110100000011111001101101011000011101010000000111011011111000010111111000110110111001111010011110010011010001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1957[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1957, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011111000001001100011110010111011110000001010101011101111001000000110101001011011110001000101000100111101100111011010111000010; 
out1958 = 128'b10101111011101101000111101111001110111000110000001110001011110000111111011110011111011001111000110101001110100010101110001111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1958[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1958, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101000101011110011010100111110000010011101010000101110001000011101110000010101010011000100001000010011000110010011001001100; 
out1959 = 128'b10100100011111100001111011000010110001111111001001111111111001101000111110010110111010010110011101000001000100100101000000101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1959[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1959, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000101100011111011100011000111010000001011010010001101111101001101110100010011011101000111000001110011101010011100100100001; 
out1960 = 128'b11111010010101100100111111001001001100110101100101001101111001100111011000110110100000100101110100110110100010111001010001001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1960[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1960, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110001111111111101111111111010111001011001100001101100100110101100011010000111001110001000011110011110110001001001101010110; 
out1961 = 128'b01000011010011100101010110110100111111000011000101000110111101111011000001001000110111001110111010101101001000000101001001001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1961[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1961, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110101010000101101010000010010110001111000101000001110010001110010111111011111111100101101011011001111011010110101001010011; 
out1962 = 128'b00100111011111010001110100000111110111101110111001000011000010100001001001100010100110010011111111111011100000001011000100101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1962[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1962, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100001110100110011001010111111111100010000000100100010101111011110100111000101100100110010111000110000110100111000101000011; 
out1963 = 128'b11111010101001001110100100011001101010011000100011110101100010111001100001110110011110110001110000001110001000111111010110100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1963[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1963, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010010000100000101001011110111100110000011000111110011010010001100011000101110001111101100111100000101111101000010001101111; 
out1964 = 128'b01110001011001001100101110110101011000101101011001101011100010100011100111110010000000010000010001100000111100100111110000100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1964[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1964, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000000100111100101001010101110000010101100101110001101000000101101101000011111111110100010101110010111000100111000000000100; 
out1965 = 128'b00111100110110001001011110011001000011010111111011100110010111110110001001011101100101000011110001010000110000011100010110010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1965[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1965, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010111111110100110111010101010100111101011011110000010111001011100001100000011011001000100101101000110100110110000101100001; 
out1966 = 128'b11100011010000111011110100100110110011000010100000100110000010101000000011101010011001111101101101111101001011001000000001010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1966[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1966, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101110010110000101100011100010101000010010101101100101010000110101111000001110110000001101110000111001000010100101101111111; 
out1967 = 128'b00000101101111100101110011000101001001111011101010010010111111001101100001010010010000100011011101010100111101111111110001110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1967[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1967, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101111011001001110011000110111110001000010010111000001100000101111101000010010010000100011101101110011100001011001010000110; 
out1968 = 128'b10111000001110000010010000100001011111010000010000111100111111010100000100011100000000010110111011010100111011011000100000111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1968[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1968, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001001101001001100101110011101101001111010011100000100000110000100101001011100011010100110101000011100100000000010100101001; 
out1969 = 128'b01001110000010011000000100000011110100101100000000010010110101111101001011010110001011111101000011100010010111010100010111011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1969[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1969, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110110111101001011100101010010111011101001101110110111100111010011001101011011010111000001000100100101111010011110101001001; 
out1970 = 128'b11100000010111010101001100010110100011011011111111011001100000010100101001111010101110110101111011001011011010101001110001000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1970[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1970, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101111111100010101001000110110010100010100000100011011010011010100111111010011010101111011111000101001111001100111110110111; 
out1971 = 128'b11100001011101011001111000110111011010100000011101011110111001110101111001011011001000001010101101101011110110000000111110011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1971[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1971, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010110001011000100010100010001001001111101110110010000011010110001101000011001011000011110110010100111100100010100000100000; 
out1972 = 128'b10011100100111100000110001111111111011011101001010100010101110111000101010100100010111011110010001100010011010000100001000111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1972[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1972, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011010001110000001011100011100011000101111100010100101111100111100110000011000001010101100110101010010110010110110000011111; 
out1973 = 128'b01101100011011110111010110110001011100100100000001101000000010001000000011010101010101001111100001001001011001010100000001000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1973[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1973, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100000100110111110110100101010010000010111010101010011000110001010000110111101111001010111011001111000100010100100111110010011; 
out1974 = 128'b11011111110001111011010000111001100010010101011000011001001100001100101011011110101011100100010001110011110100000101111000111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1974[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1974, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000111001111010110011001001010111101110101101100010011001010110011001011011010101011010010001000111010111111100010111010001; 
out1975 = 128'b00100010011011100100011000001000011001010001010110010110001101110110011110010111001000011100010100011111001000001011101110111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1975[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1975, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011111010011111011111111001010000110011000011000011101011001101001101000101101110100110000101110010011101100011111100010110010; 
out1976 = 128'b00010001111001000111000111110001011110000001110001100110000111100011010011011110101011100101100011100100001100011110110010010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1976[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1976, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010100101111101111100011100010110101101100011101111011011110111011010010111100011110111010110101011000001010100110110000011; 
out1977 = 128'b00110101010011100110110111010110011010001101100101101010100100001001111000100001100110010011001111110101111110100110110011000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1977[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1977, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011001010000100000000111110101001100110101011001001111001100011011100001100011101110011010100110111000010000110110110001010111; 
out1978 = 128'b01001100001010000000001100100101101110101000000011110101101101001001100010101010111111111100111000100111111110010110110000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1978[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1978, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010001111111010101100011111000010001010001110110100110100111111011000100000111110101000011100011101001101010010001000011100; 
out1979 = 128'b10101000000100000000100010100111001101001010000101001000011100111101101100110011011010000001111110001101100101001111111010100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1979[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1979, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100111010100010111101101001110011000001011010000001010000001001001011010001101100110100010010001100001100000110111010110001; 
out1980 = 128'b10000000010001001011001010110011011011100001011010111011000010010111000111011010000110110110101100011100110010111111010010001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1980[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1980, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000001000101011110100110011101011011100011110101111101100101100110010011110100111011001010010000010110101101010100001111110; 
out1981 = 128'b11111111111011010001001111100010111011010100011001001001010010000110111010110000101100010000011011110011001000001010001000111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1981[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1981, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011100110101001010110110001010100101110001101101110001100010110000111000100001001011011001100011100100010100010000110110000; 
out1982 = 128'b00100001100010110111011011100011100010101001101001111111110011101011000010000101001001011101101011111110000101011111001000100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1982[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1982, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001111010011111101100101010101100000001001110011110010011011001101001101111000010011001010110100100111101101010010011101111; 
out1983 = 128'b10111110001001100111011100001010110001000001100011000000010111100111010101010101100111001000010101010111001011001110100000100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1983[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1983, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100011011011001100100010000000011101111110100111100111100011101000010111010111001100000010011100010101100101111100110110111; 
out1984 = 128'b00001001011111100001011101101001101100011000011101010000101001010101011110001111000001011001100100000010010100101001100101100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1984[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1984, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010100010100110010101011000000010001100111010101111000011001001111001110001110010111000111111001100110111001000110001110000; 
out1985 = 128'b01010000000011100001110101001000001101000110100001010111110100100000001001000110001101110110010011000011100010111001010101010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1985[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1985, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100011111001101001010001101010110110011110110101001001000010010011000001000001011011011001100010011110010011001000001111010; 
out1986 = 128'b10001011000110100001110111001100101010111000111011010111001001111010101110010110100111001010101101000101111110000110101111100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1986[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1986, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011101111010110110111101110100111110010100010001110101011100010101001001100010000011110100000001100110101000010001011110111; 
out1987 = 128'b11101000100100111100011100100101010011110010001101101100001010110011001100100111000110010010011100011011001010010010010011101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1987[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1987, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010001001110101011101111010000111001000101100101000111101011010000100010111010010000101111001011111111001001001000010110011001; 
out1988 = 128'b11111100011101010001111001100010110000110010011101010010101000111101111111101011001011101011110001111100010000000100101110111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1988[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1988, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011010001011010001011000010110101010111101101110110100101100110000001101010110001000101111100000110001100011110111101100001101; 
out1989 = 128'b11001110100110100001011101110011101010110010101010010001101110001111001111111000010100011011010110001010111000100010010000000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1989[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1989, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101000000011101001110010000011111011100110000101001000100011110011011011111011111000101000001110101110011000110001010111110; 
out1990 = 128'b10100000011101010111111101001101011100101111100101101110011100101100000100010000001010001101101101110101001011000100111011101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1990[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1990, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001111001011101101110100001011001011110101111001101110010111100011101000000001001110101100001110100100000000010000110010010; 
out1991 = 128'b10001010011010101101011100110100100011010111111011110111000110101011100111011011111000101000110101110010110010111011111100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1991[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1991, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010001011111011100101010010011000111011000101100001011101000001001111011011110001110101111001010011000101001100011100101010; 
out1992 = 128'b10101101000110011010101110110010110100011011100000100011110000010101010111100010010101110001101101001001001110000111101111110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1992[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1992, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100100111011011001101001011100011010000011101011011000001000010000001100101110001100111111001011101111010101010100101000000; 
out1993 = 128'b10111110111011001101111001010010001010000010111110010100001101011011000111101001011010111011011000010100100011101111110101100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1993[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1993, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011111000000111001110011010110011111101100000100111000011111101111001101101110110111001110010100111100010111010000010111011; 
out1994 = 128'b00011101110011111101010010110111111010011111110000010001110000011011011110000111110100110100010011000111100101110000100000110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1994[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1994, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110010111100000111011111011100011100100100110000110111000101010000111011101110111100011011100011001010001010001111001000110; 
out1995 = 128'b01110101101111001010000110000000001011011110111001000000010110100111010101011101101011000111110001001100100101000111011010001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1995[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1995, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110000001110100100000100001011011011000010111010000010100111110100000110100001010000010101011010111110000110000101001010100; 
out1996 = 128'b10001010111110100100100001110010111000110111001010010010001011010011100010101100110010010111010110000001111000101011101011010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1996[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1996, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001101000011101011100111101000111000000101000110101000101100010100000110101101101111100010100010000001010010001000010101001100; 
out1997 = 128'b00100011011111010001011101011100111100000000100100110001001111111000111000000110100110001010101111111000111001100011010001110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1997[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1997, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000100001011110111000011011001111110110001011000101001110101111111100110111111011111110001101010110011110001111010001101011; 
out1998 = 128'b00110110110101000101011100111011010100011010011000111011010111110111010010011011000101000010010011100010101111011111110001001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1998[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1998, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110011111001111110100100011001010110101010101000000110111111010010100111000011000000001100000010000011010101100110001111011; 
out1999 = 128'b00110000111010010011111101000001001100101001010111100010001010000101011000111001111001011110100000011001011110100011100010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out1999[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out1999, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001011001110010100111000000010110101101001010110001001000100011001100000010101000001101000111101111100110001101110000100000; 
out2000 = 128'b10100001101110101100000011000111111000000110001110010001010111111110010111011111110011101100001001011101101010011011111111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2000[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2000, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110010110000000011000010010000111001010101000111111011110110000100111001000010100101100111001110100111101110110000101000001; 
out2001 = 128'b11100100000101111110010011110000000111000001010000000000010011110001110010011111100011011011100010000100011111101000111010011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2001[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2001, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100110111010111010100001111100000110111011010101011111111101000100111101101100000100111100110111010111001111001111000110110; 
out2002 = 128'b01101000100011110010100100011101110010110011111000110110101101011110101100000000011010011110001010111010111000000101000101111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2002[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2002, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010101000000110101100011111101110011101111110011111100110010101001100001111001000110010000001011110100011011000001010010110; 
out2003 = 128'b01010101101100110100110001011101100010110000001011011100110111011111100010101100111111001001000011111000101001000011010110110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2003[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2003, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011000011010110111101101011100010101111000101110001000110011001001000010100010111100000101000000001000111100000100110010101; 
out2004 = 128'b11000011001100110000011011100101110111110010001111101000001101000110101100000010011011011010001111011111001101001110011100101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2004[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2004, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101100111100110001101001100000100001000001000101011100000101010000010000010001100111000011111111000010101111111001111000011; 
out2005 = 128'b01111110111010011010111100001111011110000111100111110101011011110010001111101011110000010010000101000001001101011111111101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2005[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2005, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110111001111111001101110001101011011001111100100000101110101111100001111001110100010101101010100010010000111001011110100010; 
out2006 = 128'b01101110101100001011001001001101110000010011001000110100001101101100000010000000011100011110110000101011001000010011011010000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2006[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2006, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001110010101001000101000101011000100011101110101010000011101001000010110100010000110001100010111010000100110110111101001111000; 
out2007 = 128'b10000110001100101001001000111011111111100001011000100001101000010111101011101111010001001000101110001010011101011101010010101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2007[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2007, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111110011001011011110011011110001011000001110011011010111110011011100111101100001100000000111111001000001100111100100011110; 
out2008 = 128'b10100011000010110011100110110111001110011001001000001101100011101110110111110001110110001111110000110001001101111011001110100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2008[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2008, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010010100100001010101101001001100111011111010010010001100010100011001101111100011111100100011011111001011001110101011001111111; 
out2009 = 128'b10110111100110110110011011101000010111110101011011000010111110000100010101101011000111000000011111000100111110111011010100111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2009[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2009, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001111001101101011011110011011000100001110111010110010000101010001010110010000110110111110001011100111111000000100010100001; 
out2010 = 128'b00001110110000000110101100111100011000111011001111101001011011111101100110011011011100100000101110001011000111101011111101110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2010[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2010, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101110011000010011000111010110011110011010100101001011000100100100110011010111011001111000001110011101101011110000101111111; 
out2011 = 128'b11110110001110011111101110100001101011000100101111010110000010001110101001101001110011101011101110110010100101010000001110100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2011[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2011, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100100011001011000000100011111000000010111110001010011011000001101010111001100000011000111100010000110111011010101011011011; 
out2012 = 128'b00110111101000001101111110111011000000100111111101011100101110011110101100000000101100111111111111000000011111101010100111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2012[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2012, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011011100000000001100101001000110000111010111100011010000001101111101100011101111000110111111111101110011111000101000011100; 
out2013 = 128'b10001101100001111100111100010100011010100100101101011111001001011001011001001011011101001101101000110110100010111010000111110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2013[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2013, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111100000000001110000001101111100111100101101110001111011011111000000011110001000111000000100101001101000110111011101010010; 
out2014 = 128'b11011110011111001110110101011110110001111101010010110111111010101111110001111100100001100100001100000011110101010001010001110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2014[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2014, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111010000110101010010000010100010010100010011000100001101101001111111100000111101001010010001010001110000001001011101110011; 
out2015 = 128'b11010101100000010110001111011100101110110111010000100011101011010101000101101011010000110011110010111111110000001000111010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2015[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2015, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000011000010100011101101000010011001010000110011111101011011100011101011101100111100110000101011010100100100000110111011111; 
out2016 = 128'b10010010011010100011000111011000001011000111111001001001110100001011011011011110000001000101111110101010100111111110010100101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2016[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2016, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110011101001010001010000001111000101110111010000110011110001011011111010011111100111100000111011001011110100010000100010101; 
out2017 = 128'b11111000000110000110001101000001101100001100110110110010101110000101010001001100001101011101001011100010000011010011011100011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2017[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2017, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000000011011101010101001100000000100011110000110011011101001111100101111011100110110111010111001110010010111100100111011101; 
out2018 = 128'b01001001101001001101001011010111010111011001000000000001111101100001110101010000000100100101011101000110110001001111100100001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2018[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2018, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011011001010010101110110101101010111011010101110111010100110010010011111001111000010100010010011010101110001100100000101000; 
out2019 = 128'b00101010011000110000010001011010011010110001111100100011000001001110110011111101001100011100010011010001000011001110111000101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2019[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2019, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010110110100011100101000101000011110001111000011100000111111000010000101110001100011100001000011011001000110011001010000011; 
out2020 = 128'b01001111110110110110001001111100010011100011000001011111101000110000001001111111001100101101010001100011111010010010111010110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2020[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2020, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100001110011101110011011111001001011001101110111101011101001100101111111111110110111111111011010010111100011010000101000011; 
out2021 = 128'b10101100010111000101101001111011111100000110001001010110110111011101101101000000000111001010101000100100001011001110101001111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2021[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2021, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010010110110111111111011100100101101000001111000001010001110101000110001011001011100000111111011101011001001011111101011011; 
out2022 = 128'b00000111011101100011001010000100010011111110001011101010100010110001010001000001101111010110111111001000101111011011010110101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2022[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2022, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100001111111011001100000000011000001011011001010001001110100101010000111100011011000111000010110101110111100000010001100100; 
out2023 = 128'b10000111000110000000000100011001111101011111100001000001011011100101010100110110100001000000011011011110001011111110010100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2023[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2023, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010110101010110011100000010100100100110110100001011001101111011000100011111010000100110101111111001001001000101011010000100; 
out2024 = 128'b00011100100010011010010001111111111100010101001001101011001100111110111100000001110011001111111111011011101110100001100101010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2024[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2024, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101010010001010110000011100100110000001011110100011101000111110011001100011100000000101010110101011110010101010011100001110; 
out2025 = 128'b00101101101100000111000110101010001010101110000010100110001010101110010111001010110101001101111101001011011001001010101010010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2025[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2025, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111000100110001011111011000001100001101010100111101001101110000110001111110111000110001111011000111001000111001011110111100; 
out2026 = 128'b11111000111011010101001111010001010101101001100110111011001011000011100111010011001100100100001011000110110001111010010111000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2026[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2026, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001101000001010000001000001011110101101011100011101111011110101001101111100011000010100110011000100110110011010010001000111; 
out2027 = 128'b10110100100001010011010100110100111110011001100100010010001111001101100111111000010011110101111110000001011100011010010100011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2027[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2027, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110000100001010110111000111110010001110000010110111000110111111011101001001000000111001110010011000101101001111110110110110111; 
out2028 = 128'b11000101110111100111001000110001111100001110100001000111101010111001110011111111111101011000000101111111011010001110001001100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2028[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2028, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010011110001011100100101000111110110011000001110000000010001101111011000001001000001100001010111110011001000110000101001011; 
out2029 = 128'b11111111111000100000100011011001110100011111111011001010101010000001010101010010110101110001011100110101001001111010100100010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2029[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2029, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000101010001011110010101001111011111110110111101111100001010101111111010100010100100111100000011001111110010011101110100000; 
out2030 = 128'b11100100011001101111101101100100010001111010010101101011000000000000001111010011000010000000011110110110001000110100010010010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2030[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2030, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100111011101101111100101111111001011011010100001101010010011100110001101111110110111110100101001101111001111010001111011110; 
out2031 = 128'b01111110110110010111011001011111010011100001100111110110110100011010110111001111011101100010100110010101111111000110001100100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2031[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2031, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011000110100101110000010010101011110100011010100111011101111110010000100011010111101001001000010100010011011111011111111011; 
out2032 = 128'b11101010111110100100000100010000011101101110100001000100000011101010010101101001010110001010000001100110100001000010011010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2032[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2032, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011000000000011000000011100001010010001011100010001111010101111001111111010011101110101110010100010110110110101110101011000; 
out2033 = 128'b01100100000110101110111111000111100101010011011001011110000110000101111111101010101110100011110100100100001000101101011101011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2033[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2033, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100101010111010110111101110011011001011001011111001101011000011001011001010100001001011011101111111110100001100110100110101; 
out2034 = 128'b00101111110010111000001111000110010011101111001100100000000111110000111101010010100101011111101011101011011011000111010111001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2034[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2034, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110000101010100110110011001101001110101111111001110001100000110001011110000001101101101110101101010001111100110011011100001; 
out2035 = 128'b10010001110111100001101101011011101010111011101111100100001000111011011111011100000111110011110100100100011110100110110110011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2035[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2035, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111110010101100111000011000111110011000111110100011101001101000101101010001001001001000101111010110100101100101011110110010; 
out2036 = 128'b00101111101000110001111100010010010001101111101100100110110101001100001011111100001001110001100001111100100101000110100101101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2036[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2036, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101001110100000011010000000100110001101111101001100001001010011001000010110011000010100101110010111000010110111010110100110; 
out2037 = 128'b01111011011000111101000011101001101011000100100111010111110010000010100010101000110100011100110000010111100110111101100001010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2037[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2037, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000010110110100110000010001110100010001000010001001000101101010101110000001001100111011100011011000011000011001110000111101; 
out2038 = 128'b01111001010011000010001010101110110001110100110101011011001011100001111101101000110000100001011011110001111011010111010100110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2038[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2038, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100110110101010010101101110001010111011010111110001010101100111111000001010110001111011010100000011111100100110110000101101; 
out2039 = 128'b01011000001001101110111101010000110011100100011101010000111110110110010001010000101001000111010100100111000001001100101101000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2039[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2039, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110110110111001100000100000100010010111000100011010111000001111011000011010100001001011011110100111001100100110010110001111; 
out2040 = 128'b00001110111100111111001001101000111111010101111101000101001111110101110000000111000101100000010000011111001111011111010010101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2040[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2040, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110010011001100110010000101010000101001110011011001001001100100011001011001101010110001010100000001001001110000010100001111; 
out2041 = 128'b10100110111111100011001111001011110000110100110100110011001001100000000110010100111000110101010110011100011111111101010000011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2041[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2041, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001001011110010010000110000011011010001000111001101101000100100111011100111000101000010011010111010010000001000010110001001; 
out2042 = 128'b11000100111011010011101111011111001101010101110000010001010111001110110001001110000010000010100110100011101110001000111110101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2042[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2042, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111010011011000000010100010010110101011101100100111100010100101001010000100101101110111011001111110110101011100100010000101; 
out2043 = 128'b00010001011000100111010010101011000011111010000001100110101100010000100100010110000010000001000110001110011010110001110110101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2043[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2043, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110100011100001011010101110001010101010011001011010001101111010100110010011011111111000110101101111001111001110100010001010; 
out2044 = 128'b00010000000111111000101100100111010000110011101011101101001011110101101011011110110010000000010101101001110110011010001110000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2044[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2044, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001100110101101001010001011110011001001001100111110001111101111011001100010101001011101000000011001010101010111001111100101; 
out2045 = 128'b11001010110001000101101110110110111100101110110010010101110100100101110110000010000101011011011111111011000110011000010001011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2045[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2045, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100111110110011111110010111110101001111111001111000010011011110001110100001100100111101100110101110101000101011001000100100; 
out2046 = 128'b10000100110010001101011101011000111110110000000010111110101101110110101001001100111010011010110111110001110100001111100010100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2046[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2046, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000000001011100100010001011101101111011001000011110101111001010111010100111110100101000010001010110000011011100100000000110; 
out2047 = 128'b01011100011011110100000011110100010010000101010100110010110111100011101001000111011110111010110011111011000111001011010010010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2047[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2047, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010010101100000101011111010100110100110011100010100011111001111110111101010001110011011110001010011000001110000010011011010101; 
out2048 = 128'b10111001010000001101001000101001001100101001101000111011111100111011011110101111011111001100110110001001110101000010110010101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2048[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2048, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011001111011100110110001010000001001010101001011011010100001010110000101010001001010100111011010101000001000101000110011010; 
out2049 = 128'b00110010010111111000011000000111000101100001000101111111110001001100011001100001001111011110000111001100111100010101000010001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2049[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2049, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111111111000010001101011011111010011011100101101000011110010000100101111100000111001111001000101101101011010011111001110001; 
out2050 = 128'b00110000100110110000110100110011110110110101011100000110101111111100000000011010010101101010100110111010010101100110001011010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2050[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2050, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000010100011110010010110011111111101000101101011001011010010101100011111011111101010000010001001110110010111111010001111010; 
out2051 = 128'b10000110100110100100110010010001010011111110011001100100011111101101000001011000111011101101010111010010100100011111101111010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2051[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2051, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101111101010101011111010111000011000010011100011010110001000001000100111000101110101011110110000100001011100110111111001010; 
out2052 = 128'b01001001100110110001000100110100101101100110101010001100000111111111000100011101010100001110111110100011101110011010011000010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2052[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2052, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010011000000011111111100010011011100011000110011010100101001101111100010110001000100100101010110011111000111100010100010111; 
out2053 = 128'b10110111000101011011001010010111010001110000001000110001100111000000000000010100100011001111101001000000101100011011010001101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2053[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2053, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110100111101110110101111100111011000110001110111010101110100110010011100101101101100110001011001110100000001011100001000111; 
out2054 = 128'b11000100111000010010011111000100110110011100100001111101010100011000011001111101101100000000111101010000001011010101011011101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2054[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2054, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110101100000110101011000111100000110000110011111011110000100011000011101001111010011100111110110111000010010101011011101000; 
out2055 = 128'b10111011001100001100100110000111000001000100001111101101000111000010100111000100000011010111010110010011011010010001010000100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2055[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2055, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011101110101111101000010101001001111100111000000101011101110111101010000011001111010000100001011011100111010111101001100100001; 
out2056 = 128'b11011011100010100001001100100001111010001011011110000100011011011100111100111100011001010101010100100110111000110001000001011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2056[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2056, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001100110011110101100110000000100010001010010011001001101101011001110101100011101111111111010001001010010000011001011000010; 
out2057 = 128'b10101101101101111100111110111000011110101111011110011101000100110010000110100100101111100000110111010000111111010000111000100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2057[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2057, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100100000000010100100110101111001101100001100000011011111100111011111111010101010101001111101010100111000001111110000011110; 
out2058 = 128'b10000001101001111011010110011110101011111100100000101100011010011100010010000001111101110100000010101001001101011111000101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2058[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2058, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000000001011111010110110111101001101101000000000010100110111011101100100100010110011001110110011111001001010010111000111001; 
out2059 = 128'b00001000101011010101100110100000111100000111010110111001011001100010111001100011010110100101011100001010101011010100101001011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2059[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2059, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001001111110001001111110001100111000000001001100000111001011011010110100110101110000101110001001011110101100011010001011001; 
out2060 = 128'b10010101100101001001001011110010111111100111100010110011001111011100001111111000010111010110100010111100000110010100001010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2060[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2060, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110000100000110101011100111010111111000100111000111011100011100110010100100100000111100110111101111100111010011110100100001111; 
out2061 = 128'b00001110000010010000110111100111000010111111000110110011100010011000100111110000110110110001110010011010110111010111110000110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2061[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2061, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110010011010100010000100000111111101110001110011111110101010110110010000110011001000100110010001100011100100010000100001010; 
out2062 = 128'b11111001111000111001111011110000111110101100100110101100001111001000100100011001110111011110000101001011111001101111101110000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2062[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2062, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110111000110101001100101101010011111010011111011101011010101001010110111011010000110101011001101110011101001110100100001110; 
out2063 = 128'b11111001001110111000001111001011001010001110110110111010110000011011001100000000110111111110100101110110010000111010001110111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2063[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2063, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111110111001011000110111110101110001100000110000010100101110100100101001000100110101001111110110110001011111111100100011101; 
out2064 = 128'b01100100101111111110111110111000101101010000110000111010011011101101101010011011110011101110000001010111110011111001010000111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2064[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2064, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101100101100010101110010001101100001001101111000000100001010111101010000000100000100000100101110100111000000100100110001001; 
out2065 = 128'b00110011100001001000110010001110001111111100001111111011001011010110101011011101100101100100100110110011011100000000101100101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2065[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2065, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011100011001010100010111001000011010010000111011000110000110001001110100010011111110111101111111111110010111000110110000010; 
out2066 = 128'b01110110101110111000100110001000101010001001011011110000000000111111001100101010110101101110110101001111010111000010011110101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2066[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2066, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101011011101101000111001010000010111000000001000100001010001001000111011110111110100011011111011101110011011010011110011100; 
out2067 = 128'b00101101011010111010010101010100111111011001111001100100111111001011000011011011100101011101100011101000110100110001100101001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2067[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2067, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001010000100000011100011010111110001001111100100010010000111000011010111011100101110100001110100101001111011001111100010111; 
out2068 = 128'b10011011111010001100100101110100111010011101000011000110000111010111101111010000101101000010110001100000010010011001100000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2068[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2068, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110000100111011010010110101011100000011001100010111010110000011010011101000001100101101101110101010110111010000011110110100; 
out2069 = 128'b00001001010100100111100101101100010001001011010101101101010011110100010101001100101110110111111000100111001101011000000011111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2069[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2069, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111001011101011011111001000010111001001101010001110110000110110101011100110010000100111000000110000011111100100110100100011; 
out2070 = 128'b00101010011111010110010011001100001001111000110010001001110100001011101111101101101011111101011001011110011011010111001010110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2070[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2070, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111010111011110101011010001010001100111101110010101100010110110011100101000011011100011000010111111101100001001011111010011; 
out2071 = 128'b10001111100001110001110000110010110011000011110011111010001110111010001010111101110110100111100100100000110011001001011001000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2071[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2071, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000010011000100101101100001101100000101000110001110010101011101000011101000100111001010110011011100010000100100010101101100; 
out2072 = 128'b10111100101100000110111011001110111110011100001110011101110111111000110000110000000010000100011100001111110000000101000010011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2072[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2072, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001000011100011111110001010010001010000111101101000000111000101101110001100111011100101011011001000111011011001000001111100; 
out2073 = 128'b01111000001101011010100100100001111001001100011011111000110000010101000101100010110011000001001011000110101100100111101100111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2073[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2073, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010011010010010011011000101111100111010101001011100000010100110000110000010000100010001111010110101000111100110110000110100; 
out2074 = 128'b11110110101000001110100000110001110101111001111001000100101011001101101010001010110001011111011101010001000001000011011111010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2074[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2074, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110010011110101010001001010101101000101001001001011100001100100100010111101111111011010111010111000011010111101011110011111; 
out2075 = 128'b10111011100111111010111001100000110110100100011000110111001011011010011000001000110101100110110110011010000101000001000101111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2075[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2075, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010001111100110101010011111010010111110010000100111111011100011110001000011000011010000010100101100110101111100000010011011; 
out2076 = 128'b01101000000101111000001101111101110011011110110011011111110001001111001110110110000000001010100100011001101001001001001111111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2076[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2076, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010010111100011011010010011011010110110100011000000000111101000101101101110010000100001111011101011111111101100001101101111; 
out2077 = 128'b00001101011010010101111011101101111001110101111111111110100001000101100000001000110001100011101111101110101010000000100111011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2077[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2077, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000100111101111011010110100101101111110111000110110100111000001111110011010001110100011011010111111100001001100100100100100; 
out2078 = 128'b11000100000111101110000100110110110011101000011110011011100101001000100110000101011101011011101011000010111100101100001101101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2078[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2078, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111100101001111001001111011011101100110000100011100100010010101000111010000100110000011000110000100111101110001101001110111; 
out2079 = 128'b00101100111101011001101011111000100100000111111101101000101000100101111111011101001011000001100100010110010111011111001111100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2079[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2079, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001011011011100011000001010110111000111100011101000001100100001000001101000010100001110110000110000111011001101000100101111; 
out2080 = 128'b10100111111101101101011011101100000010111001000010000110000011000110110110111000101010000110001001101110010011010100000101111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2080[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2080, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010001111010100000111000000101011000111010010000010110100101010011010011000010111110111000010100100101111011101001000010000100; 
out2081 = 128'b11100011111011010111101011010010010100101101100100100010001011100001111001100010110111101110010110111110001001100100111011011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2081[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2081, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010100101100010111111011100010010001001110101100010001001011001010011100010001010110111101100101010101100100100001011110010; 
out2082 = 128'b10100000011100010111001111001011100100101100010110010011001111000011100010111100000111001000100111010101101011011101001001010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2082[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2082, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011110110111111010101110101111010001111010001110110110010010001011110111001101011100011011010000110001111110000100000111000; 
out2083 = 128'b01100101000101100001101100101000000001001000000000000100000111100110001011010100101000000010000011011101101110011111110000101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2083[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2083, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101000100111110010111101100100101010111000100000101001011111000001010001001100011000010100001000000000010111100110011110001; 
out2084 = 128'b01110110100110101011110001111101000011000010111001100010100100100110111000000111000101000000011000001101100010100101101111010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2084[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2084, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000010011101000101000000100011110101110101111001000010011001001001110000001100010110010001110111101101101100000001010000011; 
out2085 = 128'b01101001100101110111000011100001001011001011101000011010001101001010110000110000101100101000101100000001000011000010010010011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2085[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2085, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110111001000111100101001011100000100000100011001100011100010001110011000000110110010110101100100110011011111011001100111000; 
out2086 = 128'b10010001000111001001001100000100101001011010001100000100101101111110110010010100010111110111011101100101010000010110001100101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2086[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2086, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010101000111010011111110011011100100101010001110000000001011011111011110100111010001110111000010110010011011100001100111011; 
out2087 = 128'b11000111101101011000100100010010000101011001001101101000100101111101110010010110000000010111001001011100000011111011100111001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2087[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2087, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101001010101001100000101100001011100100010011000111011001101100101101011101111111000110010011100011010100010000001100100011; 
out2088 = 128'b10010011000011111100101000001100001011111010100001011010011101100100110111100010010111001100000111011001111100110101000100111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2088[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2088, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110001000100101101000001101011000100101011011000111000111011010100100011011111000110101110101110010001100011010110001110000; 
out2089 = 128'b10000100010000111100100101111000010110101110001100000000000110101101011010011010111001101010110100010011001010110111101010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2089[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2089, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110001011110001111011011001100001010001100011100000000011001101011101001010001101101100111100001010010000100000010000001011; 
out2090 = 128'b11001010111001111101100111001110011000110111100101010000110111010010111111100011110011101100000111011111110101011110011000011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2090[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2090, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011000101101001011010100100101111011001010010100101010101001001100101011111100101110111110101111010110011110010101010010111; 
out2091 = 128'b10010111101010000111001010100001000011000100100000101011000110000001101000001111000100011110010010110001101110100000111110001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2091[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2091, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000011101001100010000100010011111101111001100100001100000101010110001010100011010110011011110001100110111001001110010101001; 
out2092 = 128'b01101100011001001101101001101111111000100000101100110011001111100011110110000000001100010110100000111101010100110110101101001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2092[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2092, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110110001000110110000010111010110010100001010100111110101110000111010100101001111111010100001110010001001000001101011011010; 
out2093 = 128'b11101111011101000011111111010101010100010010011111000111111001100010110100010101111100100000100010010011111001000011110100011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2093[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2093, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100001010001010001010100010100100010001011111000111101010001111110011010000101000011101011110010010011001001011111101011000010; 
out2094 = 128'b11101001110101100010111101101000011010010001000011100001111010010100011110111111101000101010010000111111100111100101110100011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2094[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2094, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001000000100101000111010010000111000010100101000100110001100101011110010000111110000100010110110111000010001100000101111010; 
out2095 = 128'b10100111100000101100001001001010110010011010100000010101111100111001100101101000010001110010111110111101110100110001111001111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2095[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2095, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101011110101011001101111110011000100101011011100101111001111001101101110000000100111010110001000110011110100001010100101011; 
out2096 = 128'b11000100101100000110110010100011000101100111001111011001000010101111001001001010101100010100001101011011010111010010000110000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2096[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2096, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110100000100101001101011001001110111110101111110111011111000001110001001101011000010110010010000011000011111001100010011111; 
out2097 = 128'b10100111010110101010100001011011110000111000011010000101010110101101111001100011001000111100111111110111000000111100010011110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2097[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2097, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111100011000100101111101001011111110001101011110110101000001000101000111011000011110000110011011000011100010011110111011001; 
out2098 = 128'b11100101011011111011110110110010010111001101010010110101100101100110011100010101111101100001111101110111000110011010111111001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2098[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2098, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110101110001110101111100011111111101101111001110000011110010011010110111101010000010111110111101011111111000001110100110110; 
out2099 = 128'b00000101101101111101011010110101011101101010100110011001001100101111010000000110000011001100000111100111001101001000100010010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2099[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2099, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010110010000001000100000110000001111011110101011011000011000100101011001101111101011000100011000100010001110001111010110001; 
out2100 = 128'b10000000011000011111011100000111101101110110100110001111000101111100110010011010101011001111000010110000011000101000110111011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2100[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2100, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010110110000010000110111111000000010111100110101001001101010010101111101001100000110011110011110110001100111101010101100100; 
out2101 = 128'b10000100011110110101111010110011100100111101110100011101100101010000001111100011001000101111110011010111111101100010010011110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2101[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2101, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100111010110010001000100001001000000010101010010001011000100000011111101100011100101110000011110100011110110110001010010100; 
out2102 = 128'b10000100100001000101100011000011001001111000100010011111100101000110101000010001011100110001110001010010101110010010101000011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2102[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2102, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011000110010101110100000010010000110011011011000011001111000100101000101100001000010101110100111001100110100101000010100000; 
out2103 = 128'b11001100011100001000011111110110101010111101001000001000011110010001100010011000110110100000100011110110100000001110000110101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2103[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2103, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010101011100011000101110001010111011010010100001001101111111011011111000011100001011110001001011010001101101000010000100111; 
out2104 = 128'b00010001001101010011100111111100101101011000111011000111001110111101001110100001001001010010101111110101011010010110110010000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2104[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2104, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111000101101011000111111000110011111111111001010101101100101010100001011000000101100111001001000110011011010011010101101101; 
out2105 = 128'b00011101000100111101111100110101001001100101101001001100000101100111001100101000000110111111000010101010011100110110000010011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2105[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2105, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001000100011110110110100111011001111100011100111010001001011101111010101100001111001111000100000101011111011110100011010001; 
out2106 = 128'b11011011000000011000110000100011110011111011001001111010011001011100100000011001100110010010001010111110110100001010010011100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2106[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2106, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111000101000000111010001110100001101000000111010110110100111010000111101010001101101000111101111111110000010110001101011110; 
out2107 = 128'b00001000100011100000100100111001101110001000000001100001011100011010111001011100110001110000001100010100100101011110111111000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2107[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2107, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110001101110101101001101110100101100111011100011011011100111100100101011101110100001111000101110111010111000101110110100011; 
out2108 = 128'b10001100100000100010100011000001110011111100001101111111001011111001101100001111111001100101001001100011101101000100110000110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2108[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2108, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001100001101001001110001001011010000100001011101101000101001010001100101111010001010110000110010100110010000110100100100100; 
out2109 = 128'b10101010110111101001101000010011100101000011010001101100100010001111111100100011101011001001011001011111110011000010000000111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2109[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2109, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110000110101011011111000100011010000110011001010011110011110110111001101010110010000010111100011110010100111111101000110101; 
out2110 = 128'b11000110010110010101110011101110110110010110110111101001100100111010110010010010101111011001111110101000101101001110100010100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2110[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2110, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110011010111100101101111001010010100110000010101000000010000001100111100000101100000110100010101111001111101010000000100011; 
out2111 = 128'b00100100110111000010011001010011001000001011000101110110010010001000110100001011110110010001010011000001010100101000111110000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2111[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2111, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110100000010101011010100110100011110110011111011011010010010011100010001010011110111110010010101011001000001110011101000010; 
out2112 = 128'b01100010010110001110000101111110101011000000100011101001000000111001010110000010110111100111111001110111010011001110101000011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2112[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2112, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110101000100101010100111001000100101001001010010001101010000000000001100011110000011111010110101110000101101100000101001100; 
out2113 = 128'b10110000011101000111010000100111011001111001011011001110000011111001111110011110111000110001101011010110101111100101110111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2113[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2113, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111011110100011011010101010010001111100101101010100010001100011111111001010111001110010100010100110111001110000010100100101; 
out2114 = 128'b11110101111101100011101111100101000110000001100110111100101100011101001111011100111001010101010111000111010010000000000110000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2114[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2114, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011110111011011101110000011011011011010100010010011110001110111101101010011100011100001110110011110100010101100111011101000; 
out2115 = 128'b11101010101010010010001101001000001010101110100001000010111010011000000010110001000100110101001000101101011000011110010000111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2115[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2115, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110011100011101111011000111110000011010110011011010110010110100110110101011001010011110110110101101100010111001001100011100; 
out2116 = 128'b01000111101011110010011000111000110111001000000001111100100001110001011101000100100111101000111000100101101111010010111100101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2116[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2116, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010011100000001010011101110001110001010011101111001110011100000110110010010001111001111010110100100111100101001011010111000; 
out2117 = 128'b11010111100010100111100101111010001111001001110001100000100100110010011010101000001000011001110010011001100011010100010000000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2117[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2117, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001101011100010000010101100001110111110000111111001001000101101110110011011011011111100011110111010100100000001000010011001; 
out2118 = 128'b01101100001001100001010000000111110001001100011001111110010110011001111010101000111110110000100111010100000101110110011110101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2118[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2118, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101001001111010101011110101101000001001001110101011111010100001110000011100101010111111110111111011110001111111111011001111; 
out2119 = 128'b11011001110110100001010110000111001001110110000110101000010011010110101100011010010100111101101000000101101101110100010101110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2119[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2119, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001111000111100101110000100011011011100010010101111000101111000011111110110001111100111011001110010000010101010001001100011; 
out2120 = 128'b00101111000101101010010010010111101100011101000011101100100100011000011101101100011000101000101101000101101111111011111010000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2120[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2120, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100101100010000101010111101010011001011010110010000010011100010111110000111001010000110101010010000101001111011010010101110; 
out2121 = 128'b00111101011001010010011110010001101111001000111011010111110101100111010101000110001001111101011010101101010010001010111001000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2121[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2121, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000110000011110101110100101101011100010101100100110001001001000011100100011000101111101110110000010000011001010111000001100; 
out2122 = 128'b00100101010111110111010001000110110000001011011110101100110100000011100000000011010010101011000001010110110010111011101001100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2122[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2122, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000000110110110101110111010110010000100101110000010100101110000101100111010101000100010011100010110010100110001010100110011001; 
out2123 = 128'b11001001111000110101010101100010000010110101010000010011111011000010100000100110100100000011111000100111100101011101110110111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2123[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2123, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110011101011010110101100011000111001110001010000101000100111101111111101011110100000111000010011001011100010110011100000010; 
out2124 = 128'b00100000101010000001111110001000110110000110100110001000000110010110011010011011111011011111111110111011011000100100011110101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2124[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2124, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101111110101010110010110111111111110000100111110110001001110011000000001100011001011110011000011000001100101111000001001101; 
out2125 = 128'b11010110000010000101110110001110001010010000100000100010101010111001011100011010001001001111011101011000110100101001000011001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2125[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2125, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010001010101001110001001101001101011001110110101111101001010010001100011001100011100111001100010110011110001110000110011001; 
out2126 = 128'b11110110110100110001000011010000111111100010000101011100011000111010001000010100001111111100111000111110101110111100100101111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2126[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2126, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110000001010000011110100011001000010101111010001101100011110111001001100101100010111100011001000111010110100001000001001001; 
out2127 = 128'b01110100011111110000111100010110000011101011011100001010110000110011000101100100001010111110110101101100110101000000000000100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2127[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2127, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001000010100010011011110110111000011111001001111001011010101000010100101111111110100111001000110010001111110011100111001000111; 
out2128 = 128'b11111001001000100100010110010011100001111100000100111001111100110111010111110110110000011001100111111101011011010000100110100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2128[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2128, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000011110111101001001011100100111110110000111010001111010101110001000010101010111110111111001111111101001001010100101000010; 
out2129 = 128'b00101010100111000100101110000110010101001110101111001100010101010101100110000011000000111111110011001101100110110010000110111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2129[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2129, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010011010100000000010110101001100000011010110000001100100000101110110000101101010100111111011101010110010000010100101101100011; 
out2130 = 128'b01011111100011110011110001110101011010110101100001110110010110110000100011100101000101010011100011001011101011101000010000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2130[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2130, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000111000110110111100010111100001010011111001110011010011001110100001000110101001111101011111100110010001101101010010100011000; 
out2131 = 128'b11010011011111101010001111110110001001011010010000010111010011101111000100001000011001011100110101001001110101011101111110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2131[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2131, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000101000011100110011011010010001100110111001001001001111111100101001110101010001101011101010001101000001000101111101000101; 
out2132 = 128'b01111100100010010100011001101101111001111001101101101110100011001111101000111000110101111000111101011100000101000010100010000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2132[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2132, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111110111111110001110110111010001011111010110100001001101100110100101110001111001100001010010010000001110110000000010010100; 
out2133 = 128'b00011110000010001011010110011110000101100000010100001010110001110111001111111010010111011111100101011001010110001100011000110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2133[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2133, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001110000111100011000110010101111110001011111100111111001110010100010111010111101101010011001101001110101011000011100000110101; 
out2134 = 128'b10110101101101101010111010111001011001100100101111001011010000101000101001111001101100000110011001110011111011011001000001000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2134[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2134, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110010001100000110001110101001101000110100111100001101000101001100011010101111010101011011111001100011111110110101011111101; 
out2135 = 128'b00000001011010100111010010111000011111101110100011111000001111000100101001100100100001001000101001100000000100111010000110001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2135[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2135, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101111000101000100101111111100101000011010011010011001110000000110000010000011100001100101101011101000101110111001101111111; 
out2136 = 128'b01101111110110100011010000100111101000001100011101101001111101100000101100100010011010100100001000110111000100110010110010000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2136[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2136, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001011001001111010011111000000101111101111000100110001110001000101100000101010011000101011100111110111111111111110100011000; 
out2137 = 128'b00010011100000100100010000011101010100111010111100010001110111110010010001110101101111011110011011010001011000010010001101011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2137[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2137, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011101100001110110110100101011010011000000110101010000111011010001011101100111001000001110001000110001000100111110110100010; 
out2138 = 128'b10101101100001011100100010001010110110100111011011101000100001000011100000010011101011000111001001110001100000010111011010010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2138[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2138, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011101101000000110111100001110010100000110000101001001001000001111010000111000011100010111010010000011001001111100110100001; 
out2139 = 128'b00010100010011101010101001001110111111011001011001000000001110011101011111010110010110100001111110101100010110101111000101110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2139[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2139, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001010010110011000011100011000110110100011000101101011011000110011011111000110000101111011100011001011100111001101011000000; 
out2140 = 128'b00001101110100011010010100111010101011110011101011010000000110110111010011110110000110000000011100001101011000101100010001100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2140[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2140, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000110100001010000010101111001010111011111010111001101111010000001011000110101100101101001111010100110110001000001000110111; 
out2141 = 128'b01100010110010100111111101001011101110110011000100000010000001100100110101110011001110000101100100010111011100001100010001011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2141[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2141, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010111100100110010011101000011011110010110100101101111100010100110010011101110110101100110011111111101010000011011111110111; 
out2142 = 128'b00011101100010000011100101110011000001000010111101011111100010101100010110100011110010010111010011110100001101001010011111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2142[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2142, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011011011111010100010111110101010100100011010100011101100101000010010011111011111110001101111010100101011011101100011101110; 
out2143 = 128'b10011100000010101100100000100100111111000001110101011000111000101111100101101000111000011100111001111011000010011110101001101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2143[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2143, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111111010001110110010111110001110011100000111100110101011010011101011111001000111110111111111101000100000001101111111111111; 
out2144 = 128'b00000110100001100101010001010010100001010010101010010101011111100111111000110110100111010110010011111011110100011011010011100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2144[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2144, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100100011100111000100101011101000110000101110010101000001100011110110100100101000000110001000001001011110000110111101011001; 
out2145 = 128'b11010011111111010001011001101000011100011111101111000110111100010011110110110011100111001010101011110011111000000101010100110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2145[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2145, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101010001011101000011000001111001001010110010000001010110000001110110011001101011100111111100101001100110110011011010110100; 
out2146 = 128'b00110010001011011101000110000001011011111110111001100111101111010100001100100110100100010001010101111111110111100100101110011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2146[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2146, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100000110001110101110000000110100010001101101100010110101001100101111100111000001111100101110100010011100101000001101001000; 
out2147 = 128'b00010010010110011010000010110101101010111100111111001001001111011100001100100101010100100110011110111011100001000001111110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2147[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2147, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000010000100011000000010001111110010000110001011010001000011100111000110100010001001100111101010001010101001011101010000100; 
out2148 = 128'b01001110111011000110101110100100100101011111000101101001111111001000101101111001100011000000011110011000001001010001101111000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2148[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2148, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111100110101011010101000001100010011110010111110011001100010011001011001110011010111000000001100000010001111011110101001010; 
out2149 = 128'b01001100101111110100011111000100111111100001111010111101101101100011010100001000110111111110000101101111111001101101101111111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2149[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2149, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000100001000011011011110001001110000011001000000110101100100101001111110011001000111001000011101010111011111001110101100011; 
out2150 = 128'b10100101110101001111111111001110111110100001011001010010111010101100000010000011101110011001110000011010101111010110000110100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2150[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2150, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011011100101101000110001001111011111111010011101110010101011001100000000110111111010110100010011001011000000010111011110101; 
out2151 = 128'b11100011000001011011100100101110000100001111011000000001100100010000010101100100111100011111100010000110000111111111010101001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2151[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2151, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001111001011001100010001001010101001101111000110111011110110110100010101101001101111001000001000100011111000010001011110101; 
out2152 = 128'b10011111100110010011110100111001111110011101010011111111011110100000111001000101001111101111010100011000111001110001111111110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2152[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2152, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001100101101100000111010111001110100010101001011110100101001101011010101000001001001100101011010011001001101111000001111001; 
out2153 = 128'b11010110000110001000100101010010110100100000100011011101001100010101101011001110100010011100100011001011001000110101110110110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2153[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2153, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100110101110011110011111000110000100000001010100100101011011101001100101101011010111011111110100011000110001000111111100100; 
out2154 = 128'b11010101110101111010010100100000011000101000010001010001101100000100011010111101011011101000110100101100010100110110100100100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2154[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2154, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001000111111011110001101001011001010001111010110100111101010101001011110011101110100100110001000111101001001010101001011111; 
out2155 = 128'b01111011011111100001100101110010110010111000000100010011000011011011011000010011101010101110110010011111101010101000111010001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2155[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2155, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010001111001100011000000101011001110001001001100011110001100101001111001011010000100101000000101101111011101001111000010011111; 
out2156 = 128'b10101011101001000100011001001000001010100100101011000111101010101010001010110100100011101110100101100111010110110111000110101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2156[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2156, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010011010111110010100011000011000101101000010101100010001001111010011101100111001011100011001010001111010111100000000100110; 
out2157 = 128'b01011101010101011100010110001110011001001111101001011010110110000010011001011011010100111111010011001000101010100010101110100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2157[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2157, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100111110110010110100111001011111010110001110000001010001110001010000110000110011010010001101010010111101001001010101011100; 
out2158 = 128'b01010011000011100100101011111110010011010110111000101100000000010111000000100101100000101111001010000101100100101001010111000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2158[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2158, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101101010010100000110001110110000110101101110011110010010000110001010110010101111001011000111011100000000001101001111111110; 
out2159 = 128'b01010010111010111010100101110010011011111111100011000111110100001111010110001111000011000001110001111001100101101101000001010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2159[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2159, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111010101010101000001101001001100000011111011011010011110101111111011110011101001000001010010000110111010011110100010100101; 
out2160 = 128'b01001111111100001001010011101010111111101010010100010001110100000000001001010101100000011000111100010001000101110000101111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2160[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2160, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011001000100001111000110000100101111100011001110001101101110010101101010001000111000111100110010101011101100101111011011100; 
out2161 = 128'b01110100001010110010101000010011111111110110100010011110101101011011100110100011010110110001101010100100001100101001010011001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2161[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2161, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011111110011011001011001111011001110110000101110110110100000001001001100111010010101100010011100010110101100110000110000100; 
out2162 = 128'b00010110011111100100110101100000011100100000100010011111111001100011001000000110011111111001001101100101101101000000011111111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2162[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2162, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111101010111100110111010100000100011001100100010100000011111011101000100100011100101110010110110111110110011111001100001110; 
out2163 = 128'b10100001110010101101011100011011111110111001011100100100101100111100011000100111110010110111000110011000111101011001111110111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2163[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2163, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001110001011100100100010011010001100011110110011000000011101011100000001110110010111011100111101000111011001010101101010011; 
out2164 = 128'b10101001101111000011011010101000001011111110111001000110110000011101111000100010101100011011111110010001100100001111110100100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2164[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2164, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011100001011110010111101111111111011011111000101010100011111110000010000100101011101110101100101011011101101110010100101110; 
out2165 = 128'b00101100110001010010010010101110000101001010101010011000011111010100000000100011101100111000000111000101111010110110000010000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2165[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2165, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001111110101000111101001000001100111000011011111000110111110101001110111010100110111101111010100101101010001001111110000010; 
out2166 = 128'b00101000011111111111010011011010100101010010010110101110001010001000111010111001100110011000010010101101000100000010101010001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2166[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2166, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110010010010111110101010001101100110001000111110110111110011010010111101001001010110010000110111000010101010010000010101111; 
out2167 = 128'b11010101111001101100111110111101110110111111110110000110110111101111010001101001110011100110101101010111000010110011101000100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2167[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2167, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000111110010111011000011110101110011001101001001111111010001001000001110010010110101100100101010000011001000000101011010000; 
out2168 = 128'b00111000000010001101011010111111111101000111100101001001010100110010111111011100111110100111000001000110001011111001100000001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2168[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2168, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100000110011001101000100000111100001000001010101001101101110100100101110100101001100101011111011110100010111001001100110011111; 
out2169 = 128'b10001001001111001101001001111100101110010100010010110100000000100010011110101111001010100011001100001011011101100100011110100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2169[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2169, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110111110010100011000100111011100110100111001111001011101100001011100101101000011110100111010111010111011100011001010000110; 
out2170 = 128'b01101000000100010001101011001001110111010110100001101111000001010111011010111000011100101111101001011000010110011111000111000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2170[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2170, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010011000011100000101111111101111010000000010011010011110111101001111010011101100001011101101111011000100011100111100000110; 
out2171 = 128'b00110001001110001110110100101000100011111111111001100010010011011100100111111101000010111100110100110010001100101110100000111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2171[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2171, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000010101101110100011100101011110011000100000110000011011101000011100000110010000100000111000100001100000110110100011111011; 
out2172 = 128'b00010100111011110101111101101010010001001001101001011001001010100000011111000011100111111011011011111001000110010111110011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2172[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2172, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101111011001100111111100010110101111000000010000101000000000101111101110011100101100100101000101100110000110000000001000001; 
out2173 = 128'b11101110110100010001001001010001110110010100111101011000011110110101010110011001000011111101011000000100001110011011010101011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2173[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2173, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001001011001101100101100011011010010111010110101001100100001000111011001110101101011111000010100011101111000110101101011100; 
out2174 = 128'b01001011100010001101101010111100000110000111000001001011100100011110011100010100110111100100001110010011000111110111001000101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2174[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2174, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110100111110100111100000110000101001111000001101110101000000101101001111000100101101111000010101011100101100010001010111111; 
out2175 = 128'b01101101010111010010011101100101011011000001001011110001111001101010100001001110100000111100100111010111011100101000110101001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2175[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2175, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101010011100010111011101010011001011010111100000000000000010011100110011101101000111001111111000010101100000110010111001100; 
out2176 = 128'b01101100010000100110111000011111010101111000001111010010011100101010011111011101010011111110100000110100000101000100101001110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2176[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2176, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100000111011111100101001000011111110011110001101111111100010000101101011000100110011101010110001011110110110011101010001010; 
out2177 = 128'b00110011000001100110011111010010010111011000011001001010000010101010010101100100010101100101010101111000110100101011001000011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2177[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2177, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110011001011101110111111000100000101010010100100011011101111010100010111000011011101000101100110001010111100000011010010111; 
out2178 = 128'b10000111001100010011101001110011100000111000000111011101101011010111111110110000111010001000001101100110011101000000001011001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2178[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2178, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000111001000110111011110100011111010000000000000100000111001010000110110010011011100010110011001000000011000100000001101011; 
out2179 = 128'b10001101010100011001100111111110111100110011110110010011101001110011010010100001000001001111010011010000110101101011101010001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2179[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2179, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000000000100001110111111100011011001111001011010001101001101011100101001100000110011000010000010010010100111110101011111111; 
out2180 = 128'b00101111001000110010110110001110001000100111101011100011110101100010101101111001010101000010101101001100010110101001110100110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2180[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2180, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010000110000001001010110010110011111000001010011100010010011101001111000001110010000011111000101010000001001101101110001111; 
out2181 = 128'b01100111111110100100111011100001010011110111000010011101011011101111110011011000001010100100101010100100110011011000111100010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2181[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2181, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101101111110001110011100010011000010000100100100001011001010000000101111010010110101001011110110111000011000011101000001010; 
out2182 = 128'b00001101111000110100010000100001110110001001011010100000110100110110010100110101000000011111010111111101011001100100001010000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2182[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2182, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100011111000010110110011011010010010111001111000010111001000010101110101101010111110011111101111011010110010010100000010101001; 
out2183 = 128'b10001011100100110101100101011001111111010111110011001011100101010100110010101000111011100011100101110001111010011100110010000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2183[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2183, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110001101111100100000101111101110001000000111001100111111110001111100011110010011111010001000110001101000010010101001110011; 
out2184 = 128'b11001000011000100100011000010000000011011010001001001000011111010101111010110100011100001011001101011101011000110010100111011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2184[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2184, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100000111111101011000100111111000001101111110001101010110101100010010101011010000101000101001111110101000100010011110000100; 
out2185 = 128'b00001010110100101101010011000001100000101101011011001110011010100010111111011000000111100011110110100010100000011111011000010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2185[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2185, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010010010001000101000100100010100010101101101010010000001000110110000000011110101100011101110001011000011001110100100100001; 
out2186 = 128'b00011000111101110001100001010000001001100101101010010000010011000010111101001011011010001010011010000001000001101001001001010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2186[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2186, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101010010010011000010100000010111000100001001001111111100001110101101000001110110101000011010110011111101100111100110100100; 
out2187 = 128'b00011001110100010010000101100000110111100110001001110100101111100000111010010111101011100000100110010000110101010010011010000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2187[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2187, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100101011111010011110100101110000011100011000011001001010010001111100001100101111111101011001000101111101101000001100011110; 
out2188 = 128'b01100100100100001101001101100111001011100001000010101001110110010010110010011001001000000100110100000101101000001011010000100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2188[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2188, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010001010111111010000010000101011111001110001010110110010110011000111000100110101111111101111011011000010011001001010111000; 
out2189 = 128'b10110111101011110010100001001101100010001000001000111111111010101110110100011010111111011100110111110011011010111011011101000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2189[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2189, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001000010000111011001011001110111110011010110001010001011101101111000000100001010100111001000110100001011000100000111110111; 
out2190 = 128'b01110110101101111000010101110101111011101001011000110011111011100110000011101110100111011010100111010101010000100101110100001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2190[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2190, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111111001110110111100110100000101011111111001110001100110011111100001101010110111010110101111110000100111001010001100110101; 
out2191 = 128'b01011100110010000001100110110010011110011010111011010111000100111011100110110010111101000100101110110011110000001011110110100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2191[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2191, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110000010101001111101011010110000101111110100111111011011010001000100001001001100010000111001101010010110011100010100100100; 
out2192 = 128'b10100000011011110000010000010110000001000000001101111101000010001010100011110110111000101101001001000110101001101111001110110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2192[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2192, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010010110011101011010101100000101010011000100011011111010010111011001100101001101100101011000001001010010100100000001101110; 
out2193 = 128'b01111010010100100101100101010111100101010001111111110111001100010001000101101100001010100000110011011010111110001010000011111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2193[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2193, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000011101110101001110100011010001010011000011011010010011010110011111100001001010110110001011111110100101011001100110000011111; 
out2194 = 128'b11010000010100000100000101100010110000011100011101101110100010101110000110110110011001101100101000010011010100010111110001111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2194[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2194, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110110101010110010010010001001101000101100010110100100001000001111111110110101100100011110100100010101010100110010010001001; 
out2195 = 128'b11011111100101110010000100111011010000111010100000001101101010001111110000011100001011100111110011011010101001110010010101011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2195[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2195, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010010010100010100000111100111101011111110101011110111100101101001001110110101010001100011110100000100011110011000010000111; 
out2196 = 128'b11110101011101010011111101100100000010101110001101011010001010110101011001011111001001101010011010111000011110011010001001101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2196[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2196, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100001100100010110001011010011110110001001101010000000100001000000100001000110110101111011010101000000001101010100100001101; 
out2197 = 128'b01101111010100000011000101011101111101110001000111111001010100010001111100010110010110101000000100110011010000000000100110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2197[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2197, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100000000110010111001011010101110000111010010101001010011111001001100110011011100100001101100100100011110110111001100100000; 
out2198 = 128'b00100010111001000010001100000011010110010000111001001000111100100011100010001100100010010111000110010001010000001100101010010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2198[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2198, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101011100010110101010000011110011010000010111100010111010110000110011101011110001000110001101001011101101011011011101010010; 
out2199 = 128'b01111010101111111011001010000010110000001011000110100000111111110110101001101010010011110000111010111100001111101110100101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2199[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2199, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000111111110111111000010101001111010101001011011001101110010111001101110011111110001001011001000111010001010111000101011110; 
out2200 = 128'b10100011111000101010001110001001000110101000111000101011101110100110010110110010100010101001001100100001100111110101001111011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2200[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2200, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110110010010100001010100011001011011110011010101110010010111110000111100000100011111111101001001000001110101101001010101100; 
out2201 = 128'b11100110100100100010000011110111001100010101011010010110110100100100011000001100001100100011010101011010001101011100010001110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2201[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2201, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110110010110000000011110000100000101111010000111111011110011111010011101010100001100100100111110010101011010000010001010100; 
out2202 = 128'b11011001101000010011001101111011000001111010100001100010000011111101001000001011110001101011100000011000001100010110011001101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2202[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2202, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010111111011110010100011111111111001110010110101010001010101110011010100111010001001111011001011000000001010111011100000100; 
out2203 = 128'b11101101100101101111100010111100100011011001111001101001001111011000110011010010101011100101101011111101111010000101000000101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2203[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2203, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000011110111101010111101010110000011110101001001001111110110110000001010101001000010001110011110111000100010000111011000100; 
out2204 = 128'b00110110011010101111100010011001100010100010111100110100010011001111010001110101110001111111010111001000011111110110010011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2204[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2204, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110010011000111111001001111111010011111001001110110001101110111100111110110000101101101100001101111001110101000000101011011; 
out2205 = 128'b11010100000110110000001000110001110100000110101000011011110011001001011001000010001011001110001000110101111111100100110110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2205[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2205, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010000000101110010011111000000000101001000011100000010001111011100110100110110000110010000011010000011011111110010110011111; 
out2206 = 128'b11110010010101111110011001010010010001101101011010010110010010100000111000011100111110111011110110011010110101000110100100100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2206[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2206, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100110101110111111000101100001001110111110011001111011010111000101001011001111001100001101101110011101011001100111100100101; 
out2207 = 128'b00001000101110100101001110000011111011101010011101000110011110001111111110111010000001100101000001110100000100001101110111001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2207[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2207, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011000011010010010110100111000001011111001011111110000001110111100111100101011011001011010011101111111101000110101101100111; 
out2208 = 128'b01000100000011001010000010010110000111011011111001011011100010011101100100001011000110000110010010111010101011100001011011100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2208[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2208, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111110000101100100110010000100001101001100011011010011001110010101000011111110010100001101101110000010011110101010110101100110; 
out2209 = 128'b11110000100111100000100110100011110110111100000011110110000010001100101001001010001100110011111000111101000100100000001011100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2209[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2209, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000000100100000000111101111100111010001000010000010111000001001001100101111100110101110001101110000100010011100101111101010; 
out2210 = 128'b11110110011101001110100100100011101010000010011101100110010100101010101100001110001000000010101001010101100111101010110010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2210[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2210, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111110011111100001111100001100110100101001001000001100001111101001010000110110000010111010100101111111111011110101010101110; 
out2211 = 128'b11001101010110000101100111110110100101100101111011011001010111000101100101101001000001111010010011111100010010101111100001010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2211[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2211, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100001100110100101110010110010100001100000001011000100100001011000011011001111010011010000100101101111011000001100001111111110; 
out2212 = 128'b01100010000010001000110001110100100001110110110001110101001000010110011111000111000010011100111000011001100111011010010100001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2212[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2212, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010011011001110010100111100110110011000111101111001001001110101110101101100100001101110011001010110111111001001111110011110; 
out2213 = 128'b10111110010000111101110001010001010100010101011011100001000010101100100011010001110101111110010100010000010011101001011011011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2213[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2213, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110010111111111101001001101111001100110000111011110110101001101000000100000000010001010100010111101110001011010110001000100; 
out2214 = 128'b10010100101011111000100011110010001000111011100110000001000111010000010010111110110101100000001111001010110011000100110011000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2214[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2214, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111001000000010010001101010101001100011000001011010110100101000011001100001010110001001001100111010100111100000001111100100; 
out2215 = 128'b11011101000111001101110111000010001001000000011000001100011110010111000101001000101100101010110110101100111000010111111101110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2215[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2215, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011101010010111100111011011001110010010010001000001100100010011100101010001000100101000010001010000010000110011010011110011001; 
out2216 = 128'b11011010110010101000011010111000110111010000001000001110110100010011000010010101100001001001010010111100100111101110011100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2216[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2216, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010000100011110000110001100010100111001110001110110000010011000100010100100111100110000011101011010111011111111011111011111; 
out2217 = 128'b10110011011011011000111111101010000001111111010110000000110101100001011100111001110111000100111010111111001101010000001101011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2217[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2217, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110110000100111100010101100010111110101111100111100111111111100111100111101100110011100110000010111110101011111001110011101; 
out2218 = 128'b10100011110010000011010001111111110110111101001100001001001100000011110001100011101111001101100000100011001111111111101110010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2218[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2218, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110001001111001010101110101000001010011000000110011110010011011110111011110011011101001010000110001010001000001100110110101; 
out2219 = 128'b10000001000101011100110011111100111101111001100001010111111101101011100000001110111001101001011100011111001110010011011001001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2219[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2219, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111010100000111110010011001100001111110010110110100001000100100010001001000011000011101100001011100010111010001111010101010; 
out2220 = 128'b10010001001010010001010011000100000101001000101101111110000010101110101000010000011011011001110111101111001000110111110010100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2220[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2220, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110111111011000111111101011001100000111010111110010000000011001001001101010010110001000010111011011010100101100010101110110; 
out2221 = 128'b01101000001010010100100111001010001101011100001111011100011000100010110110111101111000011011001101101110101101101111101100111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2221[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2221, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101110011000101010001000100101100011100010101011111100111111111111100011100010111100001001011001011011111110111011000101001; 
out2222 = 128'b00101001100010010010100000111101011111110011110001101000010000110011110111101010010000000010001110000111100111111000100000000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2222[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2222, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000010001101011100010000010100010010100101000101111101011100001011110000010000100001110101101101100011010111010010110110110; 
out2223 = 128'b10000001000010011110000001010000110111110010100000011100010100100100101100101000001000110111110011000000010000001101111000010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2223[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2223, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011011110011011101000001010100011010000100101101111110110001100100010011011111001001011010100101110111111010010100110000101; 
out2224 = 128'b01010111101101011001101000101111011000001000010101101010111110010011111110111010101110010010110100010000101000111011101010111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2224[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2224, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111100100101010001110111010100000011110001110011011000011000110101100110010110000001111101000110111100101101101110111110110; 
out2225 = 128'b11011100010110110001110101101010100001001011001110110111000010111101111010011000110011001010100100110001000110100011001001010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2225[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2225, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110001011001100010010100100010100000001011001001101011000010011010001000010010001101011111000100001010111110100001101110111; 
out2226 = 128'b00101100110001111000011001010001110100110100100010111100010010000100110111101111111010000110101110000100011010010101111101111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2226[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2226, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100001101100000101000101011001111100100010011001011010001001101101111111100011110000010111010100011010001010011001011111101010; 
out2227 = 128'b10100000101110011101110111101000101000111001010011000000001101001100100011000101100100011101000110101011110111000010111101111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2227[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2227, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100110001110000110001111010011001000100101001100101000111010110000111000101111110001000110111111101100001011000010011101101; 
out2228 = 128'b10110110111101101001001101101000000100010101010110111100101101111101110011100000011001010111000111100000010001101001001111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2228[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2228, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101010010011001010010011101110011010001010100100110010100011001110111000100110000000100100000110100111001001100100011111000; 
out2229 = 128'b10001100100111010000101000110010101010000010111000111010111011110100100011001110010111011101110000110001111101101101001111111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2229[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2229, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000111011001010010010000100010100010100110111110101101011111101011000011100110010110011111001111000011001001110000011110111; 
out2230 = 128'b11111100111001000111010000010101010000100100011110101110010110010011111011100111001100110100100001011111011101100000110101101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2230[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2230, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110010100010011001011101100010101010011100110001111000100110110110100101010010101000110111100000110111110000001011111000000; 
out2231 = 128'b10011001100000001100101101100110111010101000001110100001111011001100001000000101010111000011100111110001010011110110011000000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2231[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2231, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000110001101010111110010000001010110001110011001001101000000000110101000001001111001000000110110101001001100101010110001000; 
out2232 = 128'b11101011010001100000001001101000100011011001111101100000100100101100000100111101100100001001111101000110111100010100001011011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2232[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2232, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100111101000000001001101010100001101100011000001101101111110001001010000000111101100011001101100000011010010110011000100110; 
out2233 = 128'b01001010011110100000010101100001111010110001011000000111010100000011111111001110111110000000000110100111100000001110010011001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2233[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2233, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101101100001110111100011111011001110111110010001110110010101111111001111000100111011001111111100011100101101010011100101110; 
out2234 = 128'b00000111110000110011000010101000000110100000110010101111000010001011001001010101010111000111111110001110010001110100101010111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2234[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2234, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111110111001010100001110001101111001000001000001000001101101011110110000101000100100100011100001010101010000001000101111011001; 
out2235 = 128'b10110101000011110110010100110011011101110101100000111001011011111111110101010100110100011000110011110001110011001101101010000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2235[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2235, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011111111000001100000110001011001011011010111111111010000001011110110011111101001011011110100011111000001010010100110100101111; 
out2236 = 128'b01000000000000110100010100010011110110000010011111000100110100000000101010001000011111101100110000001000111110100100000011001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2236[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2236, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110110101000110011101110111100000111001110101010001100100001100101001100000110010100100011010000111000010010101100101010110; 
out2237 = 128'b11011011101010111100101100111110100011101011100001000101110110010010100010000101101100100010100000001000100010111011011110100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2237[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2237, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001011101001010000101100110000110110100011100100110101101100111100101010100111101101001001011100111101010110101101011010011; 
out2238 = 128'b11110111010100111111101010111100000010101101110100100001100011001001001011001111011000000010101010101011000110111010000101001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2238[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2238, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010100011100101100000011011001100100111000111000111000001101111010111111100100001000010111000000101110100000110000000111101; 
out2239 = 128'b01001011010001011010010011001001100001010010011010011100111001110010001111010010011110110100000011010101010110010010001111001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2239[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2239, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110010000101101010110001101011011001111110010100001011001011010101000111000111101001010110001010111011111000001000100100101; 
out2240 = 128'b00111110101000000011001101101110111011011010011101111111011001000111001011010001000100000000111001100100011110100000101111001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2240[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2240, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110101010000001000000100000011000000111111010101111011001100111000111111000100101000100100010110000001001011100001111000101; 
out2241 = 128'b10010111101010100011101000100010100001000011000100011001011001010011001110011010100110011001010011101001111111000100011100110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2241[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2241, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001111010001000101000001100010111011111111011010101111111101011111011110011010110110000000100111010000011010100100111110110110; 
out2242 = 128'b11010000001100101000101101111110100100110010000111001001101000000110011101011011111101011111110100110011010110010000110011001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2242[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2242, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111010100111010111101010011100101111010100001110010111001011010011010110011001100100001100110101110001011000111001100110011; 
out2243 = 128'b00111111100111101010010001000110111011101100111111110110011101101010000011011001001110000001000001100101110011101100101101100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2243[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2243, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100010010101110100100011000100101010110110111000111110010101111111110101011101101101000110010011010000000110111100001110100000; 
out2244 = 128'b11101011001110011000010010100010111100001000111101111110110010000011000011111001010100110110000101101101111101100110110000101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2244[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2244, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000101011000110011010100001000011111110000001000100011100000001110110111110000000000110011110110011110110100000000010000100; 
out2245 = 128'b00001111111100001110111110101001010100000001101000100010110011010010110010001110001101100100110110011000001001000001111100010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2245[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2245, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001101101011110000011000001000010110111000110000001100110010011010111101110010001010000101011111111110111100001011111100110; 
out2246 = 128'b10000010100101100110101110111010011101110001011110011110010110010110110010101010100100100000011110001011010001110011111010101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2246[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2246, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001110111101110100100001111001010011011110111011001010110101110011101011111000010110011001010010011010100001000000011000100; 
out2247 = 128'b01000000101010100110011100001100011001100001110001010101000100110010011100001001000101101111001101010011101111101100010011111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2247[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2247, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100001001100101011101000110101011011100010001100001011101110111100011100011010100110100101010101000101111011111110000110100; 
out2248 = 128'b11010111011101010101110100011001111101011011010001000011101001100000110011111000100100010110010101010001100111010100100011110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2248[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2248, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100101011010001011100111100000100110001111010001111100101000111001000100011000111110000000011111111000111100101001001100000010; 
out2249 = 128'b01111101101110011111101001000010000011100010011001111111010110110010100110111111011101000001011111010101111000001001101100100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2249[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2249, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110100100011110011000101000111110001100100010011011010110100101010001001000010011111001110001111101010001010110101110011111; 
out2250 = 128'b01010101111111101011010110010100011100011001001010010101111011111110110011100100011110111001011110111001011110111011011010011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2250[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2250, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111110101010111001111010110111101011011011010010010010001010111110010111101110110110001111101101011001111100000110001100110; 
out2251 = 128'b00000010011001011101110001010110101101111000011011001110000001010010101011000001101100110100011010101000101110100111000101110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2251[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2251, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001011101001011100111100111011001001000101110000011001010011100001000000100110000001100000000001011001010011111101001001000; 
out2252 = 128'b11010111101100100011010111111000111000111100101010010001010000100111010111111111110110001010010010100101000101110001001000001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2252[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2252, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100001101100110001001001011101101100101111001110101010001001110011000100011100101111001100101001110011011011000100000100101; 
out2253 = 128'b10100000111010010100100010101010100011010001111100100010010100100011001101000011111010000001001111010010011001011011001101011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2253[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2253, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101011110110100000010010010110101000001000101010100000110100010001000100110000001100011101010101111010110000001010110101000101; 
out2254 = 128'b00100001110111110101111100111001001100011110011000001000110110011100000101100100100010011110011001001000010101100000010011010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2254[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2254, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100000101001111100001011000101101001101011100110000011101101111101001101011011100110011010111110111001101110010011000011001; 
out2255 = 128'b11100111000101111010000110001111001011000000000000111000011110110001111111101001010101111010001010001001110011011010001001010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2255[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2255, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000110100010000101000100010011010101011011110010000111110000011101001101110101011100111001000001000110100101001011100111111; 
out2256 = 128'b11000011001110011010000000001111001001101110101010100110011001000011100111101000011101110101100000110100001011101000111011111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2256[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2256, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100100101111110010111000100111110100001010110011110000011000110111110000110100001000101100000001111000100101100001000110000; 
out2257 = 128'b11110100010111011010111100001100001100110110000001110001000110011101000101010110000011110100000110000110101100011100010011111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2257[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2257, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010011111001011000111101110011101010010111010110111101111101000011011110110001111001101111010100001000011011010110000111010; 
out2258 = 128'b00111101110110110011110101111111000101000110011101101101100111001010010111000111100111101000010000110110110100101010010100000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2258[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2258, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111111100100010110110111110111010111011110100110011011110000001001000010101001110101100111010001111100010001010000011010101; 
out2259 = 128'b00100010111100111100010100111111100000001000000101101011101100101111100111100010101111100010100111000101110100001111111100101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2259[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2259, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101000001001001101001000100010000011101100011111011011111010110100110100111010010110011110011011001001101010100001111011101; 
out2260 = 128'b11101110111110000011110110011011010000010100011010100011000000011011101001000100101111000100100001110001011001011001111110010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2260[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2260, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100100100110111001100111001110001110001110001101100011000111110110101011110101011001000110100000011100111010011001100011111; 
out2261 = 128'b10110101011101101011011010000110000100101010010100110111111111111100000001010001101101001011110000001010011001001000100001011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2261[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2261, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001100110110001001011100010100100010111100010101011001001011100010101110001010011001110110111011000000101001010110111101010; 
out2262 = 128'b10011100010010111000010010100001101101001110111110101100011000001011000111011011111100011111101010111101011000000101000110010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2262[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2262, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000100101001111000100000101100100011110000101011001000110101101011010110000011100110101111000000101000100111110111010110111; 
out2263 = 128'b01100110010111100100110010100111011001110110100101110011001111100110011100001111000110010111101010001111000001110001000010011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2263[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2263, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110001010110001101101111001001011010001010110001001100000000011000001100110000111000001011000111000000100010001011001000110; 
out2264 = 128'b10111000111110111001001101011010010100001001011010101000010010100111011001101110010111100101011101100000010000110001110110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2264[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2264, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110000011011000101001010010100111001111000111000001110000011001111101000010011000000001101011001010010110100001111011000101; 
out2265 = 128'b01101000110001111101011111101001011000001101011011111000110010100011110111101111100100110110111010011101000111010001010101011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2265[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2265, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101111111000001011000101010100110101101011010101100101011000101000010010110110000000010100100001011010011010010010001001001; 
out2266 = 128'b01101011100110010101101111011011011010011111000111000101101000011111110001011101010011000010110101010000110010010011010000000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2266[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2266, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111010110011010010001110110000000011001111101100010000001101101001100100100111010001000010010011011101001010000011110100100; 
out2267 = 128'b01110110000011111010011010000011100100110101110001000001101110001111001111001100100111000001101000011100111000111111110110001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2267[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2267, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101101001010010011111010001101010100010101111110111001101110100010100110010011000110011011100001010010010111111101111110101; 
out2268 = 128'b01101101010110000000001010111010011101110101100110001011000101010001001100100101011101100111011111011110001011010001110101011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2268[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2268, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101110110010110001000111010010001110000101101011000000001011000011011111001011001110001100111010100011011010000101000010100; 
out2269 = 128'b01001010001010011011110011110110011100100110011101110101100010101011000001101010011011000110110011100101110001100100100011100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2269[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2269, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001000001110001100101000100101111000000001000101111110101000000000111110111001110100101101111011000100111100110010011111110; 
out2270 = 128'b01011010110010010101100110010000001111000011100101000001101110011100010110110111111001011100001011111111000110010001001100001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2270[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2270, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111000001010111000100000011000011100110111101100010101101001101010011001110111101011010111000101100000100010011100000111001; 
out2271 = 128'b11101101110011010011001001000111010011010110100001110000000110000010100111000001001100110001011000010010100001100001000000010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2271[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2271, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110000110110101000001000100101101011001101111111010111011010010101010000110111001001010101111100010001111011001101000001001; 
out2272 = 128'b10100110110101010001001011100001101100000100111100101000000110001010111001011001100111000010101001001011111001000000101001111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2272[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2272, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001011000001111100011001101011001011010001111111010001011101100111000111111000001011111100011110010011011101101100111101010; 
out2273 = 128'b10011111101001110111001101100010011000101010010010100111000001100100011100101100111001110000011111000110110110000000001000110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2273[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2273, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000111100000111111111011110101110101010101101011000011101000111011010011100011111110110011111100000010111011001011100110010; 
out2274 = 128'b10000001101101010111100010101001101001001000000001001010010100100111110100110110110110010100100010011101111011001100000110010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2274[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2274, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101111110000010000111010011111010110101000101101110000110100100110110101010010110111110101011101010100110100001001000100100; 
out2275 = 128'b10111110110110000111010010101111011101111000111100100101000110110000001000111110101001001000001111010111011001110001100110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2275[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2275, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000010100000110000010100000110010111110010101011100100110100101100101010111110010110010011000011111101000100110000100101011; 
out2276 = 128'b10101111111100011011001101000110001110101011111101101111000101110100110101010100110111101100101010110111001011010100110011011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2276[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2276, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110111100000001001100100101101100111101110001010110001001001010111011010000001100001110011100001001101010100001100001101010; 
out2277 = 128'b11000010000100010001001101001000100001011011101010010010001001101011010001100110011000001101001001101111101001111111011100010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2277[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2277, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100000001011001111000100111001001000000001100101000100010001111101101000100000111000111100011000111111000101101111100111111; 
out2278 = 128'b00111100010111101110011110100010010100000110010010001000001100111111010011100001101110011100100001000010100111011001101110000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2278[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2278, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111010111001110100101000110100010011111110100111111111101001001111100001111110101101111111000001010011110000001101011010011; 
out2279 = 128'b01110100010100000001001111010100001110001011001111100111011111000101000010110100101101111111001110110010000100001110100100011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2279[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2279, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110001100100101010001101101011100000000101010100110010110010101111100001111111111100100010010000110110111001010101011100100; 
out2280 = 128'b11011111001010001100101110000000111110110110010010001011100101111011101001000010110111110110000100111111011101100000111101010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2280[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2280, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110110001001001001001101111110101111010111101100110110001000010001110101011111010100101000111010101001011010001000001000100; 
out2281 = 128'b11000011100011000011101001000001110111000000000010100011001010110011001010100100000111011101101001111110101001000001000111010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2281[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2281, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011101111101010001100000001000001101100010010001000010010001011010011001111101111101000110000001101001110101000001100101101; 
out2282 = 128'b01010101100100001000101010111101000000110111111100100100110010001110011011101110000011101110011111101101110000100101000000000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2282[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2282, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010010000010000110100111011111110111001111101011111001100000001101110100101100011110000010100010010111101101000100001001000; 
out2283 = 128'b00100110011010100001001100101011011111101010101110010010000101010100001110011110001100011000111101001011110101110111000010010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2283[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2283, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011011101011101111001101111111001000000001010001010010111111000000010001011010011110100100100111010111000001101001100011000; 
out2284 = 128'b00000000100110010010010001101011000100111111001100001011011100111101010100110101100011111011100100111001111000101101111111000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2284[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2284, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111110111110111001010101101101110001100001110000010100111101100111010110010000110000010100100001111111110101110101010011110101; 
out2285 = 128'b00000000001111001100110010101011011100111110101000111011011001111101100111111010110100100101111000100111011110000011010110101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2285[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2285, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011101111010000110011010111001000110001000111110111111011100010011011110110011010000000010110101110011011010001111001100011100; 
out2286 = 128'b11000101111100001010100000010011010001110001001010010010000011110011010111010000011000001000011000011111110110001101100100000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2286[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2286, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101011100000011111001100001011010001001011010110111101101001101111100101111011000100100001111011100100010011010100000000011; 
out2287 = 128'b01100011011100001101100101000000010010111001011011000000101001011001000010001011010100111001000011101100110011110100011011000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2287[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2287, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111011010100011001010000001101100100101100110110000111001001010011001011010001001101101110100010111010011001111000100010100; 
out2288 = 128'b00000100110001110100000010111101100001000101111011101001100110011101011011100010100001011000001010011010101111001111001110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2288[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2288, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010000001110110010111110001100001000111101011011010010111011100011001000011000101000110010010101010000000010000101100101011; 
out2289 = 128'b11100000001001011001101100110010111101011101101110111100011010000001000110111101110100001010001111100000000110010100000000111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2289[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2289, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111011101100110100111101100111001111001100100100111100100111001111010010011100101010110100001101101100001000010010111011111; 
out2290 = 128'b00100000101111100001100100001011110011111101111101101011001011111000100101001011010101011111101100000111000010001101111010101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2290[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2290, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110000001101110101111100110111111000001001011101000011010000000010000001111000010101010101001000100000110011010111111111000001; 
out2291 = 128'b01110111110111110000001000000011000101010000010011011011010001000110010100110010011111000110101101111000111001011111010100010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2291[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2291, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100110110100001001110101101001001100011110000101001001010000111110010010001100110011111001101111100011110111111000000011001; 
out2292 = 128'b10111001010011111000101111000011011011111100011110010110011111000111010000110000111110100111010000000101100110110111001010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2292[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2292, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011001011101111101100101110010110101111111010000010100011010101111100011111110101010010000000101111011001101010000011001110; 
out2293 = 128'b01111010000001111010100110111111010111011010100111010001001100010000010101101101000101010110101111101111100000011000101101001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2293[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2293, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001100111011100110101010011101000001101111001101011000101110000010100100011111110001110001111001111111101011001011110011000; 
out2294 = 128'b01111010001000010010100101100111010111000010111001000101110011010000101100000011111000001101101111101111101101101010010010100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2294[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2294, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111011100101110010111100001100011110001001110001100110110011100101111011111000100000001001100011111000010100010111100000000; 
out2295 = 128'b10010011110001011010011100001001000111101011011011010100001010010000011001111100001011001101110000011100101001111010000000011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2295[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2295, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101001110100111011011101000100010111011010010011011110010000111111000001010000111111001010011010111111000011110100101100101; 
out2296 = 128'b00001111001001010000110010110100110011001111100111010010010110100101010111011110100101100011110110100110000011111010001011101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2296[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2296, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001001110001111110000010001101000010001100001011100001100101000111011010000110110111110000000010010001011000001001011101101010; 
out2297 = 128'b10010000111010110100000001111010100100011100001111010111010001010001111010101011101101110110111011101101011110000011110111001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2297[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2297, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011001110011110111010101010101000110001000010001000011101011001001010011010001110101001000011101001101101000001101111110011000; 
out2298 = 128'b01001101110001111011110101001101101101100010110010101111010011011110010111100101111101011111100001100011001101110001100111011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2298[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2298, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000010111000110011000000010100110111111011001101010010010010001101010111001111001101011000000111000100111101001001101001110; 
out2299 = 128'b11011011001101100101001101101100010011111101111011000010000111100100011110101101110110010100100000010111110000001010101011000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2299[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2299, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010101001100000110010000010110101101110011001011010101110100101111000111111100111100000011010110010110000001110101011010001; 
out2300 = 128'b01111000000011100111111001001101111111101001001000101111110001010100001101110110101001111111011100011101010010010010011001110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2300[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2300, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001011110100010001111000010110101100011111110111001001100110101000011110011110000100100111110101110101011001101101011111110; 
out2301 = 128'b01010000011111001100000001011100000000100011101000100100010110001110101001000000010000000101000010101110110010000111011110010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2301[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2301, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011010011010101110101010110010110101110111100000100100000110110001101101001110011001010101010111000001110110110011111101101; 
out2302 = 128'b00001001001110111110000011110000101100111010111101100001011000101110110111000110000000110000010101101111010010110011101000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2302[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2302, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011111000111101000101110111010111001001010000010010010010100010110101001110000110111110010010101101111100100110010110100110; 
out2303 = 128'b01100110010100100011011111001001110110001100010110001010111001010010011000001000010000000000110000110110111111000010100000000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2303[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2303, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011010001111011000101101010010010100000111001100001100000001001101110010001100000111001010101100110011011000001011101000111; 
out2304 = 128'b11101001011000111010001110101011101011011101000001001100101011111110101110111011111011101100111101101001100110001111100101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2304[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2304, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010011011101011100011101100101110100100101010011101000001000100110101010011110101010000010011100100111100111001101110100101111; 
out2305 = 128'b10000101011001101110001010101000000110111101100101101010111111111111100101110000011101111100010101001011111010111100010000111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2305[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2305, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011100001001000110100001100110111011100110001010000010110100100111100100000110101010000001110100111111101010001110011101100011; 
out2306 = 128'b10001000101111011011010000001101010100100101101000000111111101010010011011111111011100001000011001100110000010010111001001010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2306[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2306, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111000100011110010010101110001110000011111101011010000001001000000010110010101000001001111001001100100111100001100011011000; 
out2307 = 128'b01111101101010000011010100010001111011001001001100110101110001001110010110101001111000111101011011000001010010011101111110011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2307[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2307, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000101101111100000010111000111110110011011101010110010101100010101011110111110011000101100110111111010111111001110010101011; 
out2308 = 128'b01100111011011010111010010101011011111100101111111111001000111000000001001110000100001001010011110110010001101111000010001010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2308[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2308, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101001011101001010101001010101100100100010000110111000001101111100110000010111101100111110001110110001011110110111010101001; 
out2309 = 128'b11001110110110100111110101000011011100101001011111000100010011010111111001011101111100100110010001111101110010100111001010100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2309[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2309, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001001101110111111001000100101111110001000100000100110100001101111101100110011011101011100011100110101101100100010001111111; 
out2310 = 128'b00011010000000101110001111000000101100110000111110111110111110111111100000110011101101101100101010000111001000100010010110101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2310[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2310, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100110110000110001110011011010010000101011101010111010011100010001100110100000101011011001111000110011101111100000100011011; 
out2311 = 128'b11111010100110011010010101110010001101100011101000001110100000001111000000110101100110111010011111110101101010100001000011100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2311[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2311, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111001010101011100011001011010010011000101101001010010001000010010110110100010000000010001011100101111001000001101100001011; 
out2312 = 128'b10101111001011000010000001111100010010111011000111011011110011111110001010011010001100110101010111101100110011101000011010011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2312[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2312, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010011000000111010011101101110011001110010111101001011010000111000000100000010111010010010010000000101101011000001000100010; 
out2313 = 128'b00011011000001110001110001100110001111111011110101111110000010100010010001010111110010001100110010001000010011110001101001010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2313[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2313, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001101101100111000110111110110000101000100100110100011011101100001100100110110100001011111101111010111010110011101111100110; 
out2314 = 128'b10111000011111010011100010001111101111110100100011001100001101010110000110010011011111001110110001110000011010101100101100011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2314[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2314, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011010111011001011110100000100110110011110001010000110000001001000011010111101111011001001111101001110110111110100000010011111; 
out2315 = 128'b11100101011001111010011101010100011001111000110100111111010100110100011110001010011110101100100001111010010000100111110010110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2315[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2315, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100101011010010000110011110101111101011011001111101011001111010001100111110101111110100100011010110100010001011011101010010; 
out2316 = 128'b00110110101011110111101101111111101001011011000011100111101111100110101111100001001010000110110101110011011100101011000011100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2316[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2316, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001111000101011010110100100110110001000101100101101110100101110001110001010000101110010100110000100100101111101100110000111101; 
out2317 = 128'b01011010011101010101010101111001110110000001111011000000011011001110111111100001000000000000010100010100101011110011010011111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2317[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2317, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101110000111101111010010110011111001000101000011010001111110010101101010000000001100111110101000111100111100010100111111000; 
out2318 = 128'b00100100101100010100001011101011110011100111100100010000000011000101010010101100101001101111010101000001001101001101101000001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2318[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2318, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110000111001110100001110001100111001100110100011101100101010010110010101001101001110110110101011000010111100011110111001101; 
out2319 = 128'b10101001100111001000100101111000011100110001100100100110101110110101000111111011100100110101000010101011011110111101111001111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2319[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2319, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010010001000010101111101101000110010011001001010011011001001101010001110011001100101010011000101100001110110100110110010011; 
out2320 = 128'b01110000110101101010101010101111000010001100011001001011001110100110100100111001010010010110101100010011001010111010111100110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2320[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2320, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101011110000011011101001010110111110110110010111110111000101000011110001111001000000001001110100010111011101000001010010001; 
out2321 = 128'b01010011100010110001001000000110011000011011111101100010111101011011101010110111110000101100100001001001010011111110110011110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2321[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2321, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110010111001111001110110011110111010000110011011111000001010110101011011100000101100010101110010110001010100000110010011011; 
out2322 = 128'b01000111011010001101001010101101110001010111100100101111011111101100000011101000111110000111100000001001011101001100111001010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2322[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2322, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011001100111100101000111000010110111110011010100101010000111101111111110010011010011111100100011111001111111000010111110100; 
out2323 = 128'b00111101000110101111010101100111001001011011000001110111001100001101100001011000000100011000100110011011111100000000000000101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2323[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2323, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010011111010111011011101101101100110011101101000011100100000110111110000000010100000110010110011101010010001111011010000110; 
out2324 = 128'b10100101010001110101100110100010110100111100000110000110110010010001010101111010100111010000110110001010000001001001101011100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2324[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2324, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001111110011011110111111011111100000110001000110110100001101111011110011011011100011111000101100000011100110100000010110010; 
out2325 = 128'b11111011100100010100110110001000101110000001011000010101000100010001011011000011100000010100010011100100000110111001111110111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2325[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2325, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011101010110010010010110000110110110001110101011100110000011111000101110011111101001111001011011010100000100111101110110110; 
out2326 = 128'b00110110111101101011110111111011101100001011001001101110101100001001100011111111001100100000111001011110111110010111100000111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2326[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2326, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010101101011111000010111010100000001111101111110100001111111000100111111111011100101100010111101101111101000101110000001000; 
out2327 = 128'b10101101001111000000011001000000110010110100000110000110100101111110111000011111011101010111000000100100101101100010010110111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2327[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2327, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011000001001101110001100100011000110011000011000000011111100110110110001010011100011100100111100111111011001010001000000100; 
out2328 = 128'b10011001100100010001001110100101011110010110100011110101100001001110000010100011111100100000101001011110100000101100110110100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2328[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2328, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000100111111010000110110010111000001110010010001101010000011011011111011001010010101011101111110110001011111001111010101111111; 
out2329 = 128'b11110000011001100101110011010000101110111110011101110101101111100010000010111011101100111010001010101101111111010111101101011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2329[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2329, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101011110110011101011000000000010100010110000101100101010100101111011011000000001101001100000010100010110001101001010001101; 
out2330 = 128'b00100100111111001111101010111011010101110100101010101010100000100101110111000001100001010001110001000111100011110000010010101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2330[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2330, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110110100011110110100100101100111100100010110011101001010011011011111001101000010011000101010100001101010001110000101000011; 
out2331 = 128'b01011011000110101010000000000011100110001011011100011111111110011001011101000111101011011101101101110000001101011011101110000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2331[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2331, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001010000001101101001000100010101101001101101000110010111101110000010110000111110100010011001011001000001100111111010110001; 
out2332 = 128'b01110101110000001100110110110011011001000010100011110110110100001110011001111000100100011111000101101101011111000110110100101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2332[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2332, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110111010001101000001110111110010110011000110101001101110111001011110011100100001100100000111111110111101010101100011110001; 
out2333 = 128'b11001111111100111000001101001111001111001101000101101110100101011111101010110011111100011111001100011110011010001000110010011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2333[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2333, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000010001010001111101010111110010100010110001010011000011000010010110100101100100101111010001101100100010010101100111100101; 
out2334 = 128'b11010100000001110011010101000101101100001111111001010111101110101001110111001001011001111010011010000101001110011001101010000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2334[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2334, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111010011010111001011111010101101110010100001011010101000001101010001010111100011001100011010111010000010010110111011001100; 
out2335 = 128'b11011010111110011110110101001101010011001001000100111000000110001011001011001110110111110110100100101100100001001111011000000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2335[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2335, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111101110110010101111100011100010111101001100110110111001111000000011100111011000000010011010110101011010110001111001111010; 
out2336 = 128'b00111101101101101010001110100110010010000101110000110100011111111111110001001001110000010111000000001100000000111010010101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2336[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2336, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101111001110110100011001101111110000101101000011100001011110111000110101110101100110001101100010111110100100111101110010110; 
out2337 = 128'b11001010111101001011101101110001000000111111001111001111110101011010001101010100011001001001100000001101010101011000000000101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2337[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2337, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100001001101100000000101000101100111101000010001111110111101000000101000101001011100000110011000111001010101010110000101100; 
out2338 = 128'b10011010011100111000101010110011101000111110001011011111110011100000000000101110110110100100100011111001001000000010101101001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2338[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2338, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110100000100111000000010111110100010111010111001101111011001011111001100001111010001110001010100100011111101011101000110101; 
out2339 = 128'b10101001101000111010010111100001101111111101001010001101100010000101110101011100110000101100001110000110010011101101111110011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2339[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2339, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101110110101111101101010000110000101111100111101011011101011100101101111001011001010100010000111111001011000011001100100111; 
out2340 = 128'b10100010111010000000111100000011001111111000011001001001011010110100110011111101011100110010111010111000110010111001100111010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2340[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2340, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101010000111101111111010001011000001000110100011101101010001111110010011111111111011010111010110101000011001110001000110000; 
out2341 = 128'b01000101011110001011011000010100110010100001111010100001110011100011010000111010100100010101100000100110010000000000000011010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2341[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2341, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101010011010001010010101000001000101101110001111100110010010110000100110000110100000010101001010100101100000000000101000001; 
out2342 = 128'b11010001011000010000001101010010001101001111010000110010101010000100101010101011110100010101100101010010011001011100111101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2342[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2342, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010110111110000010011101100111011010100111000110111101101011000111000100100110110110010101111010001100000100010000010111000; 
out2343 = 128'b11110001011100101101001010101110110001011010101011111001010111110110110010001001010100101111010010010010111000101101110111010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2343[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2343, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111011011010100011010110100111101000111110110010000101111110100000000001001010111000111010000100100110110101001100100100101; 
out2344 = 128'b11111001100001100101001111000111100100001001111010101001100111010101011000100110010000000110101110100010111101111100110000000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2344[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2344, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011100101100000111011011010010010110001100111000101001111100010001011100000111001100100001000101010110010111110000110110111001; 
out2345 = 128'b11010101101011101011001100111101111111110110011010110010100000111011000001100101111000110100000111101100111111011000110110001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2345[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2345, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110101100001001010001111100001001100100001111011100011001111001011010111001101111110100011101110001001110100001100000000110; 
out2346 = 128'b11010010010111001111101101111011110111100010011010011101011010111000100000111010100010001110010000110100011001101100001101000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2346[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2346, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110011110001010100110110000110101101011010101111010110111011001101010101110001010011010111000101000010000100110100101100011; 
out2347 = 128'b11000110100000010010111101011010100100101000001011000000010110111010010100100101111001010000100110000010111001100111100001001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2347[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2347, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001001010101010000010000001010101001111000100001101101110000001100010010000100000101011100011101010010100001100001110101001; 
out2348 = 128'b11100110010011000001101011011101111011110011001000000110010001010101000101000010011100111111001001101001110001100000101110011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2348[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2348, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111110011011111101001101110011101110010000001101111111011101010000000000000100000000010101111111010010010000000101001001100; 
out2349 = 128'b10111000100101000001110011111110000001001000100011010100001111110111011111010011101110110101110011010000000000001011100000101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2349[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2349, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000011110110011110000101001110101100110111010100110010110000110111110101011111000010011110010010001011000100001111100101111001; 
out2350 = 128'b01011010110100111001111101101110111001110000011010110101100000001010100001110101101010010111001101010100111010010110001111010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2350[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2350, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101000110111101011011011001111011111000010000100110011111010110101000000000010001110110011111010000111001001110110000000001; 
out2351 = 128'b00000011100000101001110110101001010101110001110100000111110001110111001100011000000100101100001111011010011011011100110101110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2351[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2351, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100000111101011011111011111111110011101100110011011111100101110101101011110001000011101010110110110010111010011110001111100101; 
out2352 = 128'b00101000011101010100000001110000000110110110100011101000100011011000011101010100111111011000010101101010011110100001111010100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2352[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2352, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100010100011000100010011110111101000100011010000001000011111101001001111111011011001011010011010010110100101000001001110001; 
out2353 = 128'b10100101110000110001101010000111110110101000101001001111100001111001010110111001001111001001011111110111011111011100100111011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2353[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2353, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110010011011110010100111101100011101110010101110110001110110110110000000000100001000100001110101011000100001101101101110100; 
out2354 = 128'b00010001011110010011001011101001001001110111110100000001011000011110010000101100000110101010111111111110111011110111010111000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2354[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2354, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111100001000010110100001000111000111000100001110011000101111100001100001010000111001011101111110100001100001011010001100100; 
out2355 = 128'b11110000011001110101110111011000010110100000110101001000010001101000111001001001010110001101011101101001001101000100001101010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2355[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2355, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001000101111110111001100010011110110111011110010110001101100101101010111110011011001110010101011101101011111011000010110101; 
out2356 = 128'b00001100001101011001010000111110110000101001100011000111101000011110010001111111000110011111011101101101010001110001000000010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2356[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2356, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101000011101010101101000100010101110011011101011101011010100000111110010000011001100101001011011111001100111111111000101111; 
out2357 = 128'b01011111111100111000011111011101111001001011101110100011111000101100001001110110101101001110101000100111110001010001000011001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2357[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2357, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110111101010010001110010110001110101001010011100001010010100001110110110111010101010111001110011111001100011110011011111010; 
out2358 = 128'b11010000110100000110100111000101110000001010101010111110000000110110111111000010101001001100011010101110010100100111000010001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2358[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2358, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000111001000101100100001101000101011010000100000001111001110111111111010001011110101111000100101011110110010110011110011000; 
out2359 = 128'b00011011011011001110000101111000010101011101010001011010000010001101110101011001011111100110111100001111101101111110101100100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2359[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2359, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110000000011110100011111101100011000100000000001111010100010101110000000001101000001011100010001110100101010010110111000001; 
out2360 = 128'b01100001100100101011100101110100001001100011101100000011111010100101110010110000110101111000000010010111011100000000101011110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2360[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2360, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101001000000010100100110100001101101000100000011110100111110010110110001110101000000111000111111111000101001010111110001000; 
out2361 = 128'b01010010001101100011110000111101110101111010010110111110110111100100001110011000100011100110000001000011111101010101011101001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2361[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2361, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011011000100101001100100111100110010100101100111001011011010011011111111000010001101110111100001011001010010101100100011010; 
out2362 = 128'b01100010110010100000110101010010101001001110100100000111101000010010000001011010101000001111000001101101001010101010100011000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2362[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2362, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110010110010110010010101111010001111010010000001101000100011111100111000111000100011100110010101100011101001111101000110011; 
out2363 = 128'b11101010110101100001100001010101110111011011010111011100000001000011011000010110111100101100011111000111111010011001110010111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2363[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2363, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111111111001011100110000100110111001001010010101100011001100100001101011101010001111001010001000010111011101110111011110000; 
out2364 = 128'b00110111100001110101110100001110111000111000010011010111100000010101111010010001101011101100011001001010110011010111001111101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2364[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2364, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110011011001101111001011101011000100111010011011011011100111101111111011000100101000100000001100011111100010000111101010011111; 
out2365 = 128'b00111110001111111011101010010001100001001100111010111010010110011001000010111100011110011110011000101100110101001100010011010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2365[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2365, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110110010001110000011101111000001001101000100000101111001110111010001110011001111111010111001000110100110101010111010100011; 
out2366 = 128'b01011010111010001010100000100000001011101001010111010000010100000110100110100011101010111001100000100001110010101110000110100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2366[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2366, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011011010111101001000101011000110111100010110010010010001000100011101111111010110100100100010010000010111000000010010111010; 
out2367 = 128'b01110110011110011010100011100101001110001000000010101001000101111011010001101000011001000100010001111000010101011101010101011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2367[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2367, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001011101100110011111010010110000111001001001100001110011111011011101100001000100011100100111000011011101001010011011100001; 
out2368 = 128'b10000110100111100101100001011001011111011001110101011111011011100001101010100011111000110110001110101111011010101110101111100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2368[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2368, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111011011000101110010100101010010001111010011100011110000001000001100011101111010000110011000101111001111010100100101101010; 
out2369 = 128'b01011011011010011110000111000101101011110010010100111100111101000011011000111100100110010111110000101001110110001100001001000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2369[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2369, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000000011010001000011010011000011111000011110011100101000010101001100001001101011100010110101101001111110001111100101011011011; 
out2370 = 128'b00100010110011111011111100101010100111010001111000111001001010010000101111010000101010000001100010110101000111000000011111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2370[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2370, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000101001111110001010100110010000101001111000100010110100101000100000110101100011101101010100000000110001110000001001000111; 
out2371 = 128'b10110010100000000011101001111100100101011110011101000001111110100010111110101111011111011111010111011110111101000101000101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2371[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2371, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010100100010101010011000011000000011111111111010001001000100111001100110010001000000001011000011100011101001101110100100001; 
out2372 = 128'b10000000100010010101100010001111100011010101110000010100010010001001000001101000110111001110000111000011010111000110000011101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2372[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2372, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101101110110000010100111100001011100011011111011110000111011011110000101000010010001010010100011001110110111111000110110001; 
out2373 = 128'b01011100011000011011111010100000110011110001101001111000111101010111100101101010011011001110011110011111011110000010001110010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2373[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2373, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110000011110000111000011110100001100101111011001110001101111011001010101010101011011100010110110010000001010110100111011110; 
out2374 = 128'b11001001001110100000101101101001111000101010100101100101010100000111010110101011100110101000010111101101100010110110010110111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2374[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2374, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001010010011111110110010010000111001100011111011101010011110110110010111001111001010110100010110111001001010110100110010111111; 
out2375 = 128'b11100000100111111110111111010001010000010111011000100110010111011010010110000011101001110000100000111000011100000110010010100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2375[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2375, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000001001101110100010101000110101011111010100001110101100110011110100110000111001010101100100000110111011001011110110010011; 
out2376 = 128'b01000110000010110000101001010010000011111000011010000001110010101110111110100101011001011110011001110011000001110001001110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2376[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2376, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100000001000110001011010100011101110100010000000100000010101100111001101100001000001011110000110111100101011101100100010010; 
out2377 = 128'b11111101000010011000000011011110011011111101001001011000100001001010101111001100110010100101011001011000000001010111011101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2377[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2377, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001110111101110001010010101100010101001001111011000010011010110010101010010101110001001101000000011001111110010010100100000001; 
out2378 = 128'b11100100111101101001001100011101001011100110011110001000010100100000011011111110110010111001111010010110010011010100111100110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2378[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2378, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010011111111011011011110000000010010100101011011111111110101110100111011010001011110001100011010011110111100000101111110010; 
out2379 = 128'b10001101010101001011010001010001110101100001111101110110001100101110001011000111010100010010011101100110110101111101011001101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2379[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2379, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011000111100011010000111110010111001011110001110001100011111010000010100100100011110010110111000010000101001010000110010000; 
out2380 = 128'b01100101101100011010100000010000000011010101010100001110100101010010000000101000110011101101000001101101101011100010111101110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2380[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2380, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001001000100010001011000110011001110110110011010110010011000001101100101000001111001010101011001010100010010010101001101000101; 
out2381 = 128'b11001100001000001000110100100111111100010010110000101001111000101101000100011100010100110110100011101100101010001100111110110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2381[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2381, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101110100001111101000111101000100111010010110110101111010001010110010011100110011101001101010001010011001000000110100101110; 
out2382 = 128'b00011110000011011011001000110101010000000010111000101101011001110001111010110001110111101001110111111000001101101111110110001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2382[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2382, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110011011001000100111011110111010100101101011011111111001000100000010010111100101000110011010011001000001110100100010001111; 
out2383 = 128'b00010100110110101011010001000010011101010001011001001101011110100101010000110010000001000000110001001001110101010011111110000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2383[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2383, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010010100110001010000100001101110001111111101011101110110100010111101101001101100010000100100011011001011110110101001101001; 
out2384 = 128'b10011011001000010100011111001100101000100010111000100110000001011111010011000111000110101010000111111101010001000011110010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2384[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2384, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100100101111100110000100100010000000000010101111110101000101001010011110010001111001011101010111000000000011000101100011101; 
out2385 = 128'b00001001111001111001111100110010011110010001110111110101001001101100110000110111100001110011011000101000011110101011011111100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2385[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2385, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010011011010010011101010011001001101111111110101100000010011010110000011111110000001101010000100011110111110011101000110100; 
out2386 = 128'b11100110101100101011100100010010111101000101101110010010101100111111011111000111001110111001011000000100111110111000010111101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2386[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2386, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011001111000100001101010000010001110110010110111001110111111110001000100010001101110011110001100110100011100111101010010111; 
out2387 = 128'b00000100101010101100001010100111010010011101110110110110110010001001111111011111000000001000101000110111100101100010001001001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2387[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2387, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011010001111111110100000100101110001010101111101110110111010100000001001100111101110000010110001011100011011010101111101001; 
out2388 = 128'b00100000111010111000111101111011011001100110010011111111011111110011000111100110111111000011111101000110001011101110100100100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2388[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2388, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000100111111011001110101110110001000100101010111001101110110111100110101100100100000111100010100001000110100000111101000110011; 
out2389 = 128'b01100101011100111111111111011010011010101001110001110100011111010111010011000100000010101101111111111111011010100010011011000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2389[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2389, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011001110011010110000000111011010100000111001110101010101011100011010110101101011101001000001011101101011001001000100110111; 
out2390 = 128'b11100110110101001110000011001100111110011111011101101000100101101101111001101111010100000010001011111010000101001100101111000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2390[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2390, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000000011010010101100000001000010111100110101101101010010101111110000101010111101110111000111011110110110111110001011111100; 
out2391 = 128'b01101000111110110110010011110111010000001000000101011000001101101010101110110000010000110101111111110000101011010101100011010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2391[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2391, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101011010000000001011000110111101010010000010101100111111001100110010000100101001010001010100001010010110100111000111101110; 
out2392 = 128'b11100101100100000100000101001110101101000010101100001001110101011001111100111111111000110100111000011001010011111111101011000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2392[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2392, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111101000111001101011010110010000101000001101011100010110000100111110000011001011001110000010100111010100100110010101000011; 
out2393 = 128'b01100000010011111010010010011011000011100000000010001000100111101111011000110011010111111111101001011101011010010101010000101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2393[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2393, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000100011100111011100000110000101110011110110011000000100111101100110110000011010100111101100100011001100111011111111100000; 
out2394 = 128'b00101000100111001100001011001110111011010011011110000000011010101000010111100100111001001001011000111010001100110011010010110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2394[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2394, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101011110011000111100001001011100101101001010011001001111001100011000011010001010111110111010110101101001101100100001111110; 
out2395 = 128'b00110001110101001101000010111101000100111011110010000011111001101010011000100100101000100001011000101111000100000100100101010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2395[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2395, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001011110111000011000100011100110000111011001000110101001110111010110001100100110000100011001011000011001000110101100100000; 
out2396 = 128'b11011111011010001011001100101001010110111101110111100101001001011101011000010010100001110110011101101011110100000110010110010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2396[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2396, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100100010011001100110111001011110101010001010100101011111101010100101101000011010000111100110110101100100000001101110110011; 
out2397 = 128'b10110000000011111101100011110010000100000111101011000010101011101010001101101011010100101111110111000000100110010000111000011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2397[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2397, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011101101001010000100100100111111010010100101101011001110101001011000000110010011010100111010010010010011011000000111011100; 
out2398 = 128'b10111100011000011000111011010010100110110010110101010101110100111111000010110001011100001100011110010100111111011011001001101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2398[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2398, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100011010100111011010100001101011011011111101001100001011110000101111101001000101001100000101100011100111111111111010100010; 
out2399 = 128'b00000111010000000100010011010100111001110111100011011110001011101110010110111011100010011111100101001010000011001010101110010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2399[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2399, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111011100100101100001010000001010000111111111010110101101000111111111110100001011111101010101110101100101111010110000100011; 
out2400 = 128'b11101001011000001110111101000010110110101101011011100110000010110101011111011100101011001100001111101000110011011001001001110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2400[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2400, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001000100101010101100100111001010011101101000001010001101001011011011111011111011001011101110101100001000100100101111000010; 
out2401 = 128'b11011100100111011001101101100010010111011101011010010000011011100101100100110110111111100011100010001100101000001110011111110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2401[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2401, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000000110010110010100111000111111000000010110001011000111010001100110110011010110001010000111101101011101111000100010101001; 
out2402 = 128'b10001001100000011000010111000101010011010011111101110110101001000001000010011110101010111000000001101001001000111001100110010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2402[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2402, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000011111010100111011110011110100100011011010100010101011000011001001010011011110100001011001001110100111000100100101000100; 
out2403 = 128'b10011110011100000001000001010010011010101100001111100001101000100010010001101000110010101011110111101000111101111011110111101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2403[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2403, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011010011101000011011001000110011110000010110001010101100011111001101101010011110101101010000000110010001000100100000000100; 
out2404 = 128'b00101100010000010100000011110011010110011100110110000110001100110010010110101001101011110101111000101100010000111101101001111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2404[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2404, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110110001000001101011000011101101010011100100000111001000010010111100011000010101100111010111101110100110011100100110110101; 
out2405 = 128'b10101010110000000001101110100100001011011001110110010001001000011011100011110111100101001000100111010110000111101011000101000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2405[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2405, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010110111111011100011110110011011110011111000010111100100011101101101100100100111100010010000001001001101110100000111111100; 
out2406 = 128'b11010001110001010000000100001111111001011101100111101000100001100010011111010111011000010001011011011010110111000011010111011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2406[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2406, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100010100111000001001011101101011101110001000110011010110101010110010110100110101010010111011101000111011100011101100100100110; 
out2407 = 128'b11100000110010001011110001000000011110111001111101101000111111011001101100010010000101011001100001100001011001010010010011000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2407[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2407, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101100011000100000100011001010010000010100111011001101111101100011001011111001010001001111101101111010101001111011000100110; 
out2408 = 128'b00000101000101101010001001011010110101110100000111000100010101011010110101110110101010111000000011111100101000111000000001101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2408[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2408, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000000010101111111010100010100111101111000101001111100100111111111110001011001011100101000111111111011110100110111001000001; 
out2409 = 128'b00111000000000010010110000000100111100010010010100110100011111110100001011000110010010110110011110100111111010011101010111111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2409[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2409, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100111101000100111111101101100010011000110101011100111101010111110010000100100011111011010010100100110001110001011010110001; 
out2410 = 128'b10011101100101110111101110110111111001100100101000000010001011111011111110011101000110001011100001010011101010100000010111010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2410[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2410, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011111101010001111011001100001111001001100001001110110001100000111001111010101010001011110101001101111101000111001001001000; 
out2411 = 128'b11011110011101001101110110001011001011110001010110010111100111111111101110000101110100100010000100001110100110101101101111011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2411[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2411, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011111110100011001000010001001101000111100101000001100000111110101001011000110001000100011101110010111100100101011100010000; 
out2412 = 128'b01111110100101100000010111001101001100000000110100101011110011001000000001110001111111111100011110010011000001000100100000011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2412[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2412, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100011110100001110111100011001011010100000001101111000010000010000010101100111100001110010011000111101101101100101101111100; 
out2413 = 128'b00100001110110101100110101100100010001110011110110000101100100010111001010100110011011100100011110101101111001111100110001111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2413[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2413, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111001010000010110001000101111111111100100100000000111100111000100011101010001001100100110110001100000100100000001010001010; 
out2414 = 128'b11000111100100101010111001010100010000110001011010011110011110111000100111000010111011000101001100001111001010011001110100011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2414[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2414, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100101000100010011001001111111101101101011110010100001010011101110001011101001011000111100111100111110010111100111001000110; 
out2415 = 128'b10001000100000011111110101100000100111001010101101000001101101011111001101111001101110100111010001100101111111011011111000010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2415[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2415, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100000110001100000010011011001111111001010000010010100100100010000010111011011100011111101111011101011101101010001100101010; 
out2416 = 128'b01000011101010100100110110010111100101010101011000110011001110011001110000110101000000111010111110001100101110010101011000110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2416[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2416, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001100011101110011000001111100011001110101000000011010110011011000100110000100011011110001011000100101000001101010100110011; 
out2417 = 128'b10000110010111001000010111100100111000010101110010101111101100101101001110011011000111111100110100010100000011000001011100100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2417[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2417, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111111001000010010011110000000000110101101100011011101110011010100101000110011111000010101100100011000111110111100011101100; 
out2418 = 128'b01100011010110110100110010010111010100010011001100001000110000111110010001100000110010001011001111111010110011101100010100100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2418[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2418, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100001011101110101001000001011010000000110100110100100000101110010001110000010111000001111110010000010110101000000101101100; 
out2419 = 128'b11000011101001110110100011010110000011001100001011101010011010111001001101001101000011010110101101001010010101101110111101111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2419[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2419, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101010001011111111110011101011100011111100011001010010000111011100001001110101010110111110000011000100111100101101011101101; 
out2420 = 128'b10010011001001011110011010100001111000010100101111001010010010100101010000011100111010110001010101001010011011011011011110000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2420[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2420, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101000101100111001000100000010011011001110100100001110000011110101101001110110100100001011000110101011111110100001010000000; 
out2421 = 128'b11100101101000110101111011110001101001100100010000110000001111110000110110010100100101100101100001101111101110010010011101110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2421[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2421, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100010100100011110100101101110110010110011100001110011110010011100010000010010111001111100011011011111011100001011000100010; 
out2422 = 128'b10110000100100110110010001101011110101100101001100000101111110111101111111110111000010010001001011101111011001101011011010000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2422[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2422, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101011001010000011111010010010111001111001111110111011010000100110110010101001000001001100111111010010010011110000000101111000; 
out2423 = 128'b00101111001010010011010000100110111101011101111100111010101001100000101001100111111100000100111101000000110000111111010001010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2423[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2423, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110011000001010100010111000100010011111111011001110111000100001110001111001110111110111100100000101010001110011110110001101; 
out2424 = 128'b10100100101011010110110100111111100010111011010101001000011010011100101100111100111011010001000100011111110000000110110011000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2424[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2424, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011100110110001011000110010000101101010100111010000111101101110111001111110111100101000110010110010000110001001101101101111; 
out2425 = 128'b11001100010111000100110111110011011011100110000110000011110111000111001101100000101000010111010101001101001011010110110010011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2425[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2425, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111000000100011001010001000110111110110010011011111100110011101011011000010011001010100100010011000011110111011010010000110; 
out2426 = 128'b01011101101111110000101010011101010000011010111001001011010001011001001000111100010011100100100110101110000011111001110001011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2426[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2426, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000000110111011000010010100101000100101011010000101101110001111010100000010001000001111101010101100000001111011101010010101; 
out2427 = 128'b00110001001100000010010101110100001011111000101111101101010111011001011010000101010111101111101111010001010100101011001001110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2427[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2427, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011010011101110010000101011101011110010100111111000011111110010010011011000111101101101101110100101110010111111001011001011; 
out2428 = 128'b11001001011011000110101111101111011110011100100110100101111111011101100111110010011000111111011011111010011100101111000001111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2428[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2428, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011100001110101011001010110111111001110110000111000110011001011011110010100000110110110010111111011010110100101011101101101; 
out2429 = 128'b11000110011011010000111110111110111011100101110000111000001000110100100101001001111111011100101101010000110110100110010101101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2429[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2429, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110101101100110100010101010100100011011110111100100001100011001100111111010011000101110001010000110010001100101010010000101; 
out2430 = 128'b01110110101011000010101011001101010001000101001010100000010000101101000001011010010010011110001111101010001010100100110111101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2430[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2430, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010000010001001010000001101000010010101101110000010101011001010100010000100010010011100010100110100101101001110110110001001; 
out2431 = 128'b00110110110001011101010110001101101010010100011111101000100001000100010100101100011111100000110000101010110011010111110111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2431[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2431, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101010111101001110000110010001110000101001010110001100111101001100010010110001110101010100001100011011111000101111011100100; 
out2432 = 128'b10100010110001110100011001101011010110110001101100011111101101101010110000001100011110011011111100110010011111001001010011010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2432[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2432, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001000111001000111001001010011000110000100100100110101100100101000111101100000110110001011110100111011100110100011000011010; 
out2433 = 128'b00110110111001001010000100100111100111101100000111010000101100001011110000101011111111100101100011001110000110011111010011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2433[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2433, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000101101001001111100110001001101000111011100111100101010001011111110001101001101001100101000111011101110010001101110101011; 
out2434 = 128'b01110111010001011101110110011110000011111011000010011011111100101110001001100010101100011100101001111111011000001001101001111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2434[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2434, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101110011010100100111000011010110010011011001111101010000101100011110011000000011010000011011010111000100101111111010000110; 
out2435 = 128'b01100010001100100101100111111011000110010100010011001001010001110001100001111111001100110001110100000101001111111110010110101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2435[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2435, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110001001000101011000100100010011110100100001001001110101110000111111010011010010110001010101111101011001110000000101110010; 
out2436 = 128'b01110011011001001110110001011111010010110110011101001110011111100000101110111110111011100100111000010100010010010001110101010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2436[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2436, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100101001101001000000001010111100001110001110001010110101110111100100010110001110001110001001101001101111101001001100110000; 
out2437 = 128'b01110110110100001001001110110010101011101000100011101100001111000011001000110110110000010001101111000010010111110101000001101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2437[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2437, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101011000011001100101000100110010101110010000100000111000110011111101100010110110001101000011010110011000000001111100010000100; 
out2438 = 128'b01010010010001001000001110111100000101010110100011010000100100001110111001011100010010101001111100010000101111110100100000010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2438[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2438, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100011001011101101000011100110111100001000111001011010110001110001111100000101001110010111111111100111100010000101000101001; 
out2439 = 128'b11110010010000111010110101001000100010101010000011110000110011100100010100010110101111100110011110101100011110101100100110010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2439[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2439, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100111001000010001101010001110001110010101000000000101000110000010100001011101101010000011101101110111111100100001010101001; 
out2440 = 128'b10100111111010010111010101100101100011100110011101011110110001011001010010000010100100010011001110010001000011111100101001010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2440[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2440, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111111001101101010011101110001100110100101011001010100111001010001001001001000100100110001110101001110010100001001001011001; 
out2441 = 128'b01110111000100111011111001011110001111000000110100110110111110011011101010010111001011111000011001011101001011000000111101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2441[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2441, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001111011101010000000100000010111010000001110111011110011101001100100111101001100110011101110001001111001000010111011100111; 
out2442 = 128'b00001011011111000101011000111011010111110101001001100000011010001101000000100000110011100011100011011101100101110110110100000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2442[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2442, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110001100101000000001110011101111000100000111111010000100000110010000100011000001110000000000001011101010001001101111111111; 
out2443 = 128'b11000101010011000000001110100001101001110011110000000011001000100110010111000111000101111011011111111101101101100010001011011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2443[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2443, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111101000010000111000111001101000110100111111001101001100111110010101010010010101110100101011011100111000100101010111010001; 
out2444 = 128'b10110110011101100001110110100001011101011000011110010010010111011000011101110001011111001111010001001001101011111000000001000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2444[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2444, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110100000001111010111001010101111110010000000111110101010101000000000001101101100111111011011010010101111111000100111001110; 
out2445 = 128'b00101101101011101111100010111101000011110000100010110001001000000100001110100100010111000010100010001100001000011111001110101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2445[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2445, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101000010111000110001010011001111110011000100000000101100100010001110101001000110101010100110010011011011010011110110101110; 
out2446 = 128'b00011010111010100100101110010110100110000101000000011100010000011001001100000101100010000100000101011001011011101001010010001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2446[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2446, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101010000101001111011010100001110111110100100001011101100101011011010001001100110100100111000110011100100101100111010100100111; 
out2447 = 128'b11011010111001000011000010000101000100101001100110110011100100011011101011101000011100001000000000010101111010001101001110101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2447[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2447, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101110100101110000011101110011001010110101110011010000101011000111011101101000011010110001001001101010010100101000010010110; 
out2448 = 128'b00100010011100100100001100000011110101101001011000011110001100011110111001110100000100100100100010110100010100101100010010100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2448[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2448, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110001010000101111001011110011001000111001110110110111101011110111011001011001111011110100010110010101001101111101011001110; 
out2449 = 128'b10000010011101011000111000111100111010111101000100011100110001011100110010010000001101010011010100000001010110101011101111100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2449[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2449, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000001011101000100001111001001111111101000010000011000011110000101001111000100111001010011010000010111110100001111001110011; 
out2450 = 128'b11101001011110000111000001100111000001010110111000000000010110000111100101011101010010011001101101000001101010010100111100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2450[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2450, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011000101000001010001111101001111010111010010011011111011100011001101110010100100110011101000100011001011110011010110101001; 
out2451 = 128'b10001101110111010010100000010101111101010110110111001010010100111110001000111101001111011000000011101010001110101011010011001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2451[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2451, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011001100100010001100010101111101010101101000001010100110000110001011001000001100011110111010011001000110100100000100010111; 
out2452 = 128'b11101111111010000000110110101101000010010101000001111111001100111101111100000100101100010101010110001110011010111100110110010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2452[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2452, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000111011110100100100110011010001111011001100011100111110111001111100101000000101100110011001000011010110110010101110000100; 
out2453 = 128'b10110011110000100111011110110001000001110001011110101100101111101100110011100001111111111101110000101001000010101000001000101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2453[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2453, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000101010000110000100000011001010001011010101010101000110101101001101110000000100110000110010100000100001110001110101010101; 
out2454 = 128'b11001010110110010111100111010110001101010000110110110011110011100010101001011111100011111011001110000110101001110111111000011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2454[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2454, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110110000111101011001110111000001101101101000110101100101000011110011000000110111010011101110000011110111111010000000111000; 
out2455 = 128'b00111000011110011101010011000011100010010110111101101100101111101101101001011001000100011111111101010011000001101010110100000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2455[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2455, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011100000100000000110100010001100001110111111011100110110111110110001100110101001011001101110100111010000100111111011000110; 
out2456 = 128'b00010110111010010000001000101001110010011100101010010100010001010011010001011111111010111001010110100101110110100001001011100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2456[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2456, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001100010010100010101100100111101011010000000101111111001000111110101011100101110001000000110001011010000000101001011100001; 
out2457 = 128'b00011110111011101010000011001101110010010100100100010100010001001111001111111111110111110000100101110011010111000101001001111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2457[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2457, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101101111010110010011011100110111001011000110101110101100110001001100010110001110111111001111010111010110101101101101000010001; 
out2458 = 128'b00111001001011011011011100101110011011000110111010000010111001000001101001000101010100011100110011011101011011011111101011111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2458[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2458, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001101010100100101100000101110100001000101111001101010000100100101101101111111010011010111001111000110001001111001111001001; 
out2459 = 128'b00001011010011100101110010001110100000000100100101011001010111101011010100011110000110010100111000101011001010110100110000011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2459[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2459, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110110010000011010011110010111000000111100101101001001000110101111010010000001111010111001010100000110010101001101011011000; 
out2460 = 128'b11110001111101010010101010110001101000100111011011101111100111100100100101001110100001111101111111111111110100001110100001111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2460[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2460, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111011111001000010101100000001101010011011010101111001101100001101111100111111001111010010010010001001001100110000100111110; 
out2461 = 128'b00011001111000110011100111100110100010010110001100000101000000110010111010000010101011000010111101110010011101110011001111110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2461[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2461, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111001011010000111010000110000000111001011011111010100100000110100001101110111010000001010100001001010010011101001101010001; 
out2462 = 128'b01111100110101110101000011100111011011100001101101011000010111010111001101010011001100111111011101010001111100110010010100101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2462[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2462, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001110010011111011011101001011010110101110110010001100110101111111111110001100011101100110001010011011100011111000010000101; 
out2463 = 128'b00101001010000100100000010101000010100101000000111001010011101111110100010111110101001001110010010000100111011010001010101010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2463[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2463, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100110110010101011110100010000110010010011000100010100101000001111001000100111101111010101100101110101000001010010110001011; 
out2464 = 128'b01110101110010011011011010000011101110000001111010110000001101000100011010000110000100010101100011110100101101100111010010111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2464[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2464, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111101010010100111010001010000110111001010100110101110011000010101110110101000100011001001100101101001100101111011011010111; 
out2465 = 128'b11110100000000001100111110101111100110001011110010011011010010000001100000101111100011110000101010011011011000001111011000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2465[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2465, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110011001110110101101000111110001010010100101111111101011001101000111101110011101000011000100100011001100111100111000110010; 
out2466 = 128'b01100100000010011011011110001001101010101100101101100011001001111001000101101110010111000001010000110110110100101111010000000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2466[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2466, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000101001011000011110111001100010101101100110011111111011111110000111011101111101100000100101000110111011111000011000000001; 
out2467 = 128'b10100100100101111111000100000110111111000101001000010110101011110011100100000111001011101011101101100001100000000110110111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2467[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2467, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000101011011010010100011010101100111110011100100011101010101011101011000010010000111101111111101111110010100100101001001101; 
out2468 = 128'b01011100101011100011000110001110011111101010100000101110110101100001000011111110010100000001011001110011100000000100110010111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2468[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2468, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011110111101010100010000010101111010001111111000010111111011011000001100101010100010101001000001000101110100111101101111000; 
out2469 = 128'b11100110011110010000100100100011100010001100100101011101001011011001001011100010011001011011010100000011001010001011100111100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2469[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2469, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001111110101010100110010001011011100110001011101001000001110010110011001011100111100001100111010001101001000100110110100100001; 
out2470 = 128'b11101111101101111011111010101101110001001011101110000001011100011111100100101111001100100101010010011000001000100110000110000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2470[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2470, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111001111111100001100011111111111010010100001100100010111111111110111111011101001000011000100110010101010011101001101010110; 
out2471 = 128'b00010001111110100011001101101010001111101000010111110001111010010011101011110101110001101011011001101011100110100011100011101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2471[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2471, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101010010011101010010010101101110110011000101100110100110110010000110101010110011100101111001000110010011110010100101010111; 
out2472 = 128'b10101101001101100000001100111111111011101001011001000011000111000111111100011100000111010011111001001101010010100111010101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2472[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2472, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101010000101010100011001001001110010010100111101010111000011000011110011011010001011111110100010001111111010010111001010110010; 
out2473 = 128'b01011110011100110100101011001001001001111101001000000001111010100000100011111111011011111000110010011101101001010100001100100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2473[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2473, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100010101011011011000011110110010010101001011100101110010010000101111000101101010100110001001000010000110101001101111001000; 
out2474 = 128'b11001011111100010110011110110011011110101010011000011111111101011101011011011011000011111100010111010010000011110101101110001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2474[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2474, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001110011011100110010000110100101010111001011111110011001111000011101111100100101001000011101110010010011111100011001001100; 
out2475 = 128'b11011011011110000011011001010111110011010110110110111001110000000111001010110001001101010111110111101100111000010001000000000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2475[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2475, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100111010110010101001001110111000001010001000101100100110110100010101011111011110110001010111011110110111000011001101011010; 
out2476 = 128'b10110011110010101110100001010101101111011110000010101100001011010100011100000110010000101100010100101111100100001111010110000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2476[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2476, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101101011101111110111110010001000011011011111000010010100001110101000010001001010111001001011101100001011110000011011110011110; 
out2477 = 128'b00011110100011011011000101010000011001111111110011111001111001001001000001100000011110110100110101011111100011101001010110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2477[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2477, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110011000111101000100101011101101010011011110111000100011100010100100010001010000001001110000101101000010010110100110001101; 
out2478 = 128'b11001001000011001011111011111000111110100101000111001001011000010100001011000111001001101111010100111001111001100110101000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2478[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2478, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010000111001100001011111010111100000000101011100101001010100111100011001011110011010011010101101110101000000111011010100110; 
out2479 = 128'b00001110000010010000110100001001011010100101110110100110011000011000100110110011101000101001110011101000010111001100111111111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2479[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2479, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011000010011001101000111000000011000010110000100010000001010111001010101000110100011000110110000011110110111110100000001101; 
out2480 = 128'b11110111001000011011011000001100101100011000001111000101000000000000110011110011101011011110111101111101100001000111010100010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2480[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2480, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110100010001010010100100110011101111111100011011011100100101011111100010111110110100001011001101111000001010001010011010000; 
out2481 = 128'b11001001101000000111010110000111010111110000011101001000100000101010110010100110111100100100101101010101000110001101000001011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2481[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2481, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110001111110001101011101110001101101111100111100111011111100011011110100011100100001100011110011111110000011101010111101001; 
out2482 = 128'b01010110011010001111101010111011100110111100011101101110110011110111001011100110011001010011001101110110001011001000110101000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2482[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2482, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010001100000110100001100010110011111010000001011110011011111011111110001100100100110011001110111000000001001010101001101011; 
out2483 = 128'b10010110000111011000010010010111001011101001011000010100001100000110110010111000100111101011101110101101011010110011100111000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2483[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2483, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011010111111001100110101001110100101111110000000101011001010101101100110100010111111010000010011001101001110000010101000011; 
out2484 = 128'b00001110101110000100100001110111111101011100111000110010110110010100100000110100000000111111111010011111111001100010001011110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2484[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2484, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111111111011100000001001010101011101010110001001100000110111100010011111101110110001001000101010111000111100011100010100001; 
out2485 = 128'b01011100110010100100101010010100011110101011110011101001001111001001000101000001110111110111111100111000000010110100011111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2485[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2485, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111110010100010101001100011001101110101110000011100001110100000111110001100111001100001100000000101011101101001001011000000; 
out2486 = 128'b01000110000001101101110011001100111101010111001111000001011100111100101010010111110010011110111100100101010110100011110001000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2486[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2486, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111100001100010011011100010000110110110001101111111011110010000110101101000101000011011100101000111110100011010100010101111; 
out2487 = 128'b01000101111101001011100111110001110101011100000000100100111010100101111111011001111001011111100000101011111110010100001001100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2487[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2487, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100010101110011100100110000100000000101111101000000000010011000100110001100010111111100111111001001110001111110110000100111011; 
out2488 = 128'b00001010111111011111000101000001010111011011110000011101010010000010011100110011101111100101111011101011011110010011110101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2488[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2488, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010011010100010111011101111101100101011010100010100100100001110001001100011100110110110101100110100001110011001011111010111; 
out2489 = 128'b11111001011111010111111111000011010111010101000001101010100110010001001110100010111100010111100100100111111100101100111101110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2489[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2489, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001011110101101110101001100000001000101011001101101110110000010011011011000110100011011011000011101001000111000000101101011; 
out2490 = 128'b10111100000110001111101010101101000010101001001110111010010010100110011011000110110110110110001100000111111101111010101110001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2490[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2490, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011111010011001100001011110010100110111000111000111000011001101101100000001110110001011111101110111101100100000101100000101; 
out2491 = 128'b00111011101001110000100100101001100010101011011010000001111111001111000110010100101110010111111001100001110000110001111001011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2491[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2491, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011110000011110111010110000001111001010100001101000001001001000001100000110111001100000001001011110100111110111011010010010; 
out2492 = 128'b00100000011001101000001110001010011000111101110001110101110010111101000000000010111010001010110010010100001101010011011100010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2492[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2492, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100101110000001100011100000100001111010111011101000101011010111010010101100001001100000011000100001110010110100000111111001; 
out2493 = 128'b00101111010111011111000100110011010011000010100010011101100111111000010100010110101001001000111000110101100101000001101001100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2493[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2493, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000100000110101000100010101100110010001111001001011100100111111000001111100011101101001001000100001001110100111110100011111; 
out2494 = 128'b11010011111101100111011111101010011101101101011001000111010101111110101111110110111111101111101110010011111010110100000001010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2494[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2494, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111010000011111100111111011000000110111100111001010100010111110011000010101011011100110000001001010010110110100101001100010; 
out2495 = 128'b00010111010001000010001011011111111011000000101000101111010000011100001111100010000111001100110001100111000101010110001111100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2495[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2495, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010111011011111010111000011100010111010001011100000111010001011111000011011000100001000011111110000101101011010101101011100; 
out2496 = 128'b11100100011000011101100110110000101000100110001001101000110011111011010011111111111001100111010111101000001101001111101010000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2496[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2496, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000010111111110000101010001111001101011110000001000011111101110101111010110010011010001000100110011111011000100010001001010; 
out2497 = 128'b11010101110101101111000010000001101010000011111001000010001010100111111001101111010001101110111000101110000111000011001010010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2497[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2497, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110101100100011011100010110000011010010011100010001001011110111001110111110110101110001101000000101011111000100000000100011; 
out2498 = 128'b10001100111000111001011010001010010000110111110010110001111100001001111000011110110001010011101011100111010011000001101100010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2498[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2498, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010010100111011110100010101010010011100111001010001011100011100100011000111111000100100011010000010000001000001101011001010; 
out2499 = 128'b01011010010110101001011000100000011001101111110101101101000011101010100100010011101101010001111111011000001101010111110111110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2499[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2499, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001001001010111100011101111000101001110010011001011010101010110010110001000101101110010101100011111000101101001110111100101; 
out2500 = 128'b10000111111010110101101101011001101010101011100111011001111000100101010111101110111101010000011111010111100000100000111000010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2500[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2500, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001011101101101011011011111011101011001000110001100110010100101101110101011101000000011011000101110100001100111111101100111; 
out2501 = 128'b10010001110101001001111110010001111100100100000111000110000101011100111000111100001101010110010000101101001010111001110010011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2501[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2501, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111111010010110100110011100110001010100110110010110010011101011100101101001111001101010111101010001110101100100001101001001; 
out2502 = 128'b10100111101111100110010100100001000001101110010101110111100101010000001110010010101110101100100100011001110110110100100000011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2502[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2502, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001011001010001101101011101101010010001011011100110110000101011011110001000101001010010001100000011000111110110001100001111; 
out2503 = 128'b11010001001101110111111010011111101001010011000110000100000101011100100111111011010000100100110111011000101111111101010100000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2503[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2503, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001010111010000111000010010000101111101110001110100001111001101111110110110010000011010011011100110010101100100100010101101; 
out2504 = 128'b10011011001100011110010100011110001000111011011011010110010111011111110110001111000011111111111100011000100110010100101111100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2504[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2504, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111101010001000101101001010011100001111010000001100011101100110101000001100010011111110000011010010011000010110111010110110; 
out2505 = 128'b10101000100100101100100101000110001001100010001111011000010011001111001110001000000111011100001010111110001010101011111000101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2505[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2505, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101101110010101011100111111001101010011111111100001111101000001100111100011110000111000001110100010110100011101011001101111; 
out2506 = 128'b00000001000001111100101101100111011010101011000010010010011000010000011000000001010011000100001000111101001001100101000101110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2506[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2506, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010100111110011111011110010111000111001111110110100101000011101110010101110010000000110100110010101100100001101011000111010; 
out2507 = 128'b01100011010000010000011010010101000111010001100110010000111100001111100011110001011001110111101001101100111001001011111111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2507[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2507, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001000100111101111110000110100101101001000100011010110110111100001110000010100001101010100101101010110110100000001001011111; 
out2508 = 128'b01101001110110001010001011100110001110011011111101001001011111001010000000110000000111001010100010011101011110001100111011101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2508[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2508, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111001001111011010000000110011110001110111011100110100101011110111000011000110111010111101001001111000101011011101100110010; 
out2509 = 128'b11010111011001000011101000101001111001111010011101001110010111001011000110010100100110100101100010111100001111000001001100101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2509[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2509, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010011100100000001101100001110111010100010101101010011010011100110111010110010010000001011101100010100011010001000000000101; 
out2510 = 128'b01010101000001001001110110101000101011101001101101010010111011001000001011110000000100111101111010111010010100010100011011000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2510[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2510, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110000010000101010011111100100101010101111010101011000000111001101011110001010000101001101110011111001100111100011010001100; 
out2511 = 128'b01101001010101111000100011100001001111101110101011000000001110011111001001100010011111011110100101010011010111101001011101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2511[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2511, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001011110111101111010011101101111111011011010011111110011101011000100011001110010101111000000111110101000001001100101110110; 
out2512 = 128'b01111100001110011000010000011111000110001010011000000111011111000100101010011001000111100101011110000110001001111010101110110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2512[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2512, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000011001011000001101110000001010010111011111000010001011100100101111011011001100111000110110010111010111111010010101001100; 
out2513 = 128'b10011010001011001011111110101100010100110101101101000001001001110011101001111110100111000010001101111000010000000100101111011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2513[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2513, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100110111100011001110111010000000110000110001100011000100101110001010011000010001110110110110111110101000111010100001010010; 
out2514 = 128'b11110010010010000100100010001100100111011001101110010101001000000000111010000101101100010101101001100110100100101111101111010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2514[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2514, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011001010001001000110000001110001010011010100000010011110001011010010110100100011011100010000010000110100001101101110100111; 
out2515 = 128'b11010011101000101000101000001110100110000101010001001100011001000100011111000111010010011100000110111111110101011011111110001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2515[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2515, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000001000111011010000000011100110100010110101001110100110111100111100001111010000110110101010110110010000100000011100011001; 
out2516 = 128'b11110001100001011000100011100100100000010011010101110010111000010011011011111100111111011011101011110000100001000011100100100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2516[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2516, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110110101010101111101100110000100111011100011101101100111100101010111111011111101010010011000001000100110110100101101011010; 
out2517 = 128'b00111001101101101011011100001101110100010001110110011011000000001111111001010001111100010111101101010001111000001011010010001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2517[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2517, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001010101111110001100100010000000110011011010110111010010011010100101000100111100010100101000011011011101001010010111001000; 
out2518 = 128'b10011100111110110001001101110101110110110000111110110000001001111111011000110001101001101000111011010010100011111111010000100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2518[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2518, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101011011101010111000000010111001110000000001001000000010100110101100111111011011100101110000011000100101110110001100100111; 
out2519 = 128'b10101010110011001100000111100000110110111100111100000011110011010101110111110000100010010100110010000010001110000111010100010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2519[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2519, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010101110111001110101110101000010000101000111011001010000101111000000110111101011110111001000000101110011101001110010011011; 
out2520 = 128'b11100110001010111111111100111111101010010001000110011011011101000011111100011111000100011100001010001010001011100101110100101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2520[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2520, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100110011100010100100110100011110011100011110000000001000000100000010011101001101010011100000010001100010011100101010000011; 
out2521 = 128'b10001010101010011011101101001110011010101100100101000000110100111101100001001110000100101101110000101101110111011000110000011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2521[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2521, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111010011011110101100110111100011010101010101111101110100011100010001010001101110100000000110001001111100100001100100101101; 
out2522 = 128'b01011111000111000100111111100011100000110011111111100011110100001111001100100100111010000100010011000110110001111001111000101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2522[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2522, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111001111000111011001001011110011101100100101000101110100100011001000011111110001011001010011110001101010110101111011110011; 
out2523 = 128'b00101001101001101010000110011001000111001000101000111100000011101101111011110111001010010100010001111100111101010011000011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2523[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2523, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101110111110111101001111100011111000011101000110001010110001111011101011101000011000101000111011010110010010111000001001101; 
out2524 = 128'b10111010111011101101011111110001001010110100101000100110100100001010110000101111111000011011011110011011010011110111101010100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2524[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2524, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101110010111000000101101111001011101010000110011001010001101000100000001101011110010000011110001100001001000101010010010011; 
out2525 = 128'b11110010010110010111000010100110011011101100011111110101010110110001001010001100111011110000010100011100111000000000000011011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2525[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2525, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011010001010010110110111100000000101011100111001011000001111010001001101100010001111001110001011010001100101111101001110111; 
out2526 = 128'b00101001100000110100001101110110000100111000000010000010111010001101101010100110010010101011011011001110000100111111011001000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2526[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2526, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011010101011100001110111110001101110011010110010001011101000100100100000111010100111110111000000111010111111000001010011010; 
out2527 = 128'b10011001111100110101011110001100101111110000110011100101110100000001011111111011111100000010111111010010001101110001001100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2527[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2527, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011100010110000100001111110111011111111010101101100100100110010110111000000101001010111011111001110110001100001100111010000; 
out2528 = 128'b10000000111110000100110101000001000000010000101011111010011100100011000100111111110001011000000100000011111101011110000000010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2528[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2528, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111001010100111110111011000110101100100100101011100100010010111011110101110001001011100100101001110110010100000110001011000; 
out2529 = 128'b11010111011100010010010010101000010000101010101111101001000010000110010000001011101001011011101111110100101100100111000000110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2529[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2529, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010000000100111011011010000000100111111101111001011010101110101000100011000110100000111011011110110100011110111011000000010; 
out2530 = 128'b01000011000011111110111111101010111010011001111111011111101110101010011110010011010000100010101011110110101110001111011110100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2530[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2530, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011111001111000111011111010100010001110100111010001011000111010100011001101010101100000111111110000000000100110010011101011; 
out2531 = 128'b11101111110000010010110101110111110100100110011101111010000000000000010010111100101101001101000111011100000110001001010010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2531[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2531, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100011001010010110100101000000000011000010001001110000000111110001101010000101011000101100101000100000011110011101101001101; 
out2532 = 128'b00011100101010110001110111111101100100110110001101100011101011001001100100111101110101111010111100100100101110101111100010001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2532[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2532, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001010110011010010011111100101000100110110101100011111100010100101111111111001001010000101111100001010000001100001000110101; 
out2533 = 128'b01101111110111101111100010111010001110100111101111101011010100001010001011110010000100101101100101000011000001010001010000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2533[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2533, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111001101110001111000001100010111110000110111010110110011010010111110110110010001011101000101100101101110000100001101100100; 
out2534 = 128'b01101001000111010101000101001010111111101100100101000001101101110110001101000001111001110111101100101010011011011101110101000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2534[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2534, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111101011001001000011000010110110011010011100101110011001001001011100110011110100111000100010101101000011110010111000111101; 
out2535 = 128'b01001001100000110000110101010011101010111110000011111000001100010101110111000000100000000110110010100000011010101101111010110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2535[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2535, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111110010000110000110100001011101011010001100111011100100111101000111011110001001111111111101010100011110010001001010100100000; 
out2536 = 128'b00100000110101110001010100111101111101011010100111110111010111100010100000100010110101010000110110001101001110100100101010001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2536[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2536, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000111001100111100111111000100110001110101110110111100110011101100011011011000000010011001000101110001101101000011101101101; 
out2537 = 128'b01101110111110011011100111111010110110111011111111100000110010111100010010010010110110100111010011011101101000000011000000110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2537[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2537, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011010101010100101110101000000010010100010000100010100010011001001000100101110010101001011111101101101100001011100110000111; 
out2538 = 128'b11010001111110010010110011110000000110110100100011000110000100101000110101100100101001100000110011011101100101001111010010000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2538[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2538, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111101011000011010100111110111111100001100011011000011110101001101100001111011111011011101110000000010101111011111111111101; 
out2539 = 128'b10101110110001101001000001010010000010101000001111011011010011001110100001110010111110001111000011111111010000001000011001110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2539[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2539, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101111010010000001111111100001100000000110010100101110000110000101110110110011001010001010101011011100111100101000100111010; 
out2540 = 128'b11011000001101101001100010000101011110000110010011110010100011000011010010010001001011110111101001011110011110100000100000010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2540[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2540, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001111110000110111000101001010110100001100100111110010110111001011010000110111000101111111001011010000001101111001010101000000; 
out2541 = 128'b00000100110001000101100010011100000111110001010110011101111111000000000110010010111110100010010101001101011011000111110111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2541[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2541, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101001110110010110101011000110110001101101100111011111001000110111010010010101010000100110011101101010110101011110100111110; 
out2542 = 128'b00100010001100111010011101111010000001000010110111101111011001100100111101010110000000101101111111111011111100100111001000011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2542[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2542, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110010001000101001110011111011101101011110111001010001010010000110010111011100000010010011000011000011101000110001011010110; 
out2543 = 128'b01100011110101111101010000111010110010101110111111100111001010001100000000110001100111101101101010100110110110001000010100000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2543[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2543, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100010110001011111111010110111011111010000110111100110001110001000010010110011010011110101100001010000010001001110001110110; 
out2544 = 128'b11001101000011101011111011001011110111011000101001100100010000001110101010111010011000111010000111100100010010000011000011011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2544[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2544, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011001011100100100010110100000100100100110100101000110111110100001100010100100011101101001001011111011000111100000001000011; 
out2545 = 128'b01000010101100001111111011101111011100100011101000110101011000110011011100100001011101110101011111101011011101001011000010101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2545[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2545, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111000010010000101000000010110110101000000011110000000001010001001111101111000011100011101001000111110010001110100011101001; 
out2546 = 128'b10110101100000100010001100010111110000011001100100011110011111101110101000010000100100010001010100111011101010001010111101000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2546[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2546, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111100110100101010111011110101011000101101100110010101100101010100001011010110100111111000001101000100101001000101111100111; 
out2547 = 128'b00100011000110110011101111010010101101110011110010000101100001001101011110111111000011001010010110010010100100001011011111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2547[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2547, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101010000101000010010100011010000011011111100000111100100010100010110101100101111010100111010111000000100111011100101111010011; 
out2548 = 128'b01000011001111110001011101111000111101101110001011010000101000100111100111101000111110100001011011011101000000100000001111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2548[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2548, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001100010111110000000111001011010011000110001011101100011001010000001010011100101010100010001000011001100000010000001100000; 
out2549 = 128'b00000100100111001001110010101110100010111100111111000001000010000110101010100111100001000110100001010001100111100101100100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2549[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2549, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111000010100010010101100011001111101010100111101110110100011001101010010110011001010011101000001111001101100001100001001011; 
out2550 = 128'b10110011010001100011000101110100101101000011010010010100010000101101101100110111001100111101000011111101111111101110111010010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2550[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2550, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110010100000010000011101011110010011010010000001001111011001001010011010000000100110101011100001101111011010000011001110000; 
out2551 = 128'b01100011011111010001000001111000000011100000000010101001001011110010111010000010110001000111000110100110001010001011010000100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2551[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2551, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000010111010010111110010110000110101001010000100001010010101101001000001011010110001010111010110000101111011010101001001010; 
out2552 = 128'b00010110110001010101100001110010101001101010000101000011001101010001111100101100010110100111000111000001011101011011110111101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2552[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2552, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010001100111010110100111010101100100100010110110111110100011000010100000101000000010000111000010101011010111101100001000100; 
out2553 = 128'b10011110000001001111110011010011010111111101011110000011101110011111110000111100011111101010011010100001001011101100011001011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2553[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2553, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111111110100111101000111100011100101100100001011110110110011001011000010001011011011000100111001000111010101101001011100100; 
out2554 = 128'b10101100100000110001100100010101111011100001011001100010111010110100011010011101100011101000111001011000111110101001101110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2554[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2554, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100111011000000010101101000100011101101011000100011101100010111011110000111101100000010101010000111000001010111110000111001; 
out2555 = 128'b01011111001101100100010001001101001011010101101111101110100111011011010111001010010010100101101000001000110101110111011100000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2555[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2555, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010110001001100100011110010000110111001000101011111011101000111010111011100111111100011111010011011011000011101111001001101; 
out2556 = 128'b01001101110000011010101101011101011110101111000111110010000001011100010100001000100011111011011110101101000100100011011011011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2556[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2556, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010101100000111101111000111011110010001000100101101001100011110101111100000101110011100010100000111111100101111111001101110; 
out2557 = 128'b01001000011010110110010100101001011101001101110001100111101001111011001010010000000111100011100101101110110101010000100010000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2557[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2557, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111001000011100011010101010111000101101011110000001100000101110000010000100001000010010111101011111100110100001010100111110; 
out2558 = 128'b01101100000001101001100001000110000111001100110001101110101110101000010010101111100000101100000111000010010001001101111001010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2558[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2558, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101101001001111010100110101001110110101111100110111101000111010100101111111010100111001101011010001000000010010001011111110; 
out2559 = 128'b10101001100001010110100100011001100011010101011100110100011101100101000111100101100100001111110001110111100011100011100000111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2559[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2559, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110100000101110011111001000101001001111001000111110101100100010011010010011111100101110101001101001000101100000010111110111; 
out2560 = 128'b01111110100110001111111101101101010000001000111111011010111000101111101000111111011000111001001101000100011001101001011010100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2560[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2560, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110111111001011010000110001000000101110110000000111100100100001111010000100000001000010100001011010000011101111110010111101; 
out2561 = 128'b00110101100100111110100000001000111011001100101101001101100011011110110111100000101111111100001101011010011110101100110111110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2561[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2561, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011010110000000110111100011001111101001110110000011010110001001010101000011110101010010010111101010111100001111101001000101001; 
out2562 = 128'b01001011001011000010010100011111010111101100000100101110110000010001110001110110110100100010100011101000010011011011100010100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2562[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2562, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011000110100100100101101000110111111001000101110001001001011000100101111111100011000000111010110110100110010100111110000000; 
out2563 = 128'b01011100011101011100001000100001001100101100010010010111111110110100000100011001110110011010110101100111001000011011100001101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2563[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2563, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111011110011110010000000110001011000000001100001010111110011111101111010000100010101001011011110010110010011111101001111111; 
out2564 = 128'b01010010111100100011111111010011101000001100100110110100011100011010101000101011101001111001101101011000111010101011011001001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2564[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2564, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010100011110110001111010101101111011110101110011010100100100000001001010100111111000110010010010100000100111001100100111000; 
out2565 = 128'b10011100100001010101100111101101101110000110101110010011110111110100101110101011010011110000010001111001000000000000001100011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2565[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2565, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000101100011111000011010000000001111010001100101000110010010110111010000110011100011000010101101010111111001111011001110101; 
out2566 = 128'b01000100111111011101100110110110000000110111101110101011010111110101100000010010101100010111011101010110100110011100011001011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2566[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2566, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100010000100010011011000001000111110100111100010100111101101111010111010101011110100010000000101010001101011011000110010000; 
out2567 = 128'b01001110110111011011110001001111000100101110000000011010001000101110011010001111110010110101001000110000001101011000010111000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2567[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2567, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000000010010100010010011001011100111001011101000000010100000001000000000001010000101011000100100000000011001111011100100001; 
out2568 = 128'b01011000011110010010101100000111111111000011110010100000000010101011110011110111111110010110011011011011110100011111110011001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2568[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2568, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001110111110001010101000010110010100111100001100011101100100101100110110101110001100111101011111101001100110100100000110101; 
out2569 = 128'b11001000010101101001011001111001110001000110011101101001100111101101010110101100110101101101110101000001011011000011101010110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2569[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2569, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100001100010011001010101010100000111011001010111111111110101100001010001001011100010000100010011010010011100101110010000001; 
out2570 = 128'b10001111011111101110111110111111000000100000011110000110100111111010000111011000001001001100111110011001110111101101000111100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2570[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2570, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011101010101000000100010000101010111001000110100011000011110101001111000010110100011001100000000100001100000110111101101001; 
out2571 = 128'b01110111111101100110010000111110101100111110010111101110110111001000010000010000010100001010110011001100110110111111011011101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2571[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2571, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010111110110010011110101111110101010110101010000000101101011010011000000111010011101111111001100011011000001110110111011010; 
out2572 = 128'b00000110011100011111110011001101100111011011111000110111001111100111111111001001101001010011111111001110011011011010001000011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2572[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2572, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011000100011100000000110001100100110101010111000010010110111100011110111100111100101010001010011011100011100000111111000101; 
out2573 = 128'b10000100110101100101010100110110011001010010101110001100110001011000010000011010111011010000110111010010010110110010101100000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2573[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2573, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011001101001111001111000101001101110010011111110011001000101010001111001101100111110110000011110010101111110111000111000110; 
out2574 = 128'b01010010011010010100111011111101111001111001001011000111100101000000111110101100001110010110100011110001110100001010101000001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2574[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2574, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101011111010111000001001001101101000100101101111011110100100010011011101101010111110100010000001010110000100001010111101010; 
out2575 = 128'b10101101111101000111011001011101111011011100111111101100100001110001010100101010001101100111101100100011100011010110010100001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2575[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2575, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100100101000011010110010011111100111100011000010010000001100001100111001011000000100000110101010110000001101101100001111011; 
out2576 = 128'b00000101010001000100011011100111111010000000011111010110010010110111100101101011000010111001000010101101110001011110001100100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2576[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2576, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101111001111010100101010110011010101101000000001011001000101011001110010010111001010110011000110100010100110101000000111101; 
out2577 = 128'b00011101001100000100100010010000001010011111110000011101011001110010000010011010101100000111010011110011111110101010001011001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2577[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2577, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101010110100100101011001010110000101100110000010100000100100110010110111100100110000010111101011100110111000000010110100001; 
out2578 = 128'b11000010010110001011001000101011110001001110111111010100100101100011010011001010001001010110111011001110100001001111111111101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2578[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2578, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011000101010011010000111001010100001110111110110101000000000110110111100000111111111000111100100001101100011010110011011001; 
out2579 = 128'b11001001000110001011110001011110010111000011100100101011100001010000001111110010011010001101110011000101111011001101010000010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2579[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2579, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100011111000100110110011010101000000000011011010011100100001000001100011011011000010111010111000000011101000010110110000010; 
out2580 = 128'b00011001100010100001111011100010011110011101100011100010101100110100010100011011111000011011101000110011011101110100011011100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2580[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2580, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000111010010111111101101000110011001101100001010001101001001001010011001001111111101111001101010000110110011000001111011101001; 
out2581 = 128'b01111001101110011111011101001101010000100010001001111001001001101110101010000110001100011001111110101101110111010110100111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2581[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2581, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001001110001000111110001100001111110010100001000101110100101100010000111000111001011010100011100111001100101111000001000010; 
out2582 = 128'b01010100000100010100111000010001111011101111101000000001000011000000111101100110000000000011011111110010011001010010111111100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2582[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2582, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111000110011010110101100110100100101110101100101101001100010100111000000011100100000001011011111000011010000000000001000011001; 
out2583 = 128'b01111110101001100010111010011111110000011100000111111000000000001101001111100111000100110010111010100111011000111011100111110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2583[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2583, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010100111001111101010001101001110000001100011101101110001011001110110000110110110100001100110110100101010000000101101000000; 
out2584 = 128'b00001010110000100010001111111000101101100100001100001100011011100000101100010011100101110101011110001010110000001111011011110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2584[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2584, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111110111110001111111001010110000001100101011000111110000101101010011010001010010000111111110011010000110100000101101101001; 
out2585 = 128'b00001101111100101100001111100100110111100001011001001001011001111100111000001111010011101101100100110111100110101110101100010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2585[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2585, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100110000000101100101000110001000110010001000001011110011110001011001110001000001001011001110010011000101111000000001100011; 
out2586 = 128'b01001110000101011101011000100111011010111010110010111111111110110100110010100010110110000111100111001100010001110110111000110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2586[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2586, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111001111011111011000101000011100101111100110111011010001010000000111100111001011111100101010110100100001001111010111101001; 
out2587 = 128'b00010001110011110000110001010101111000010111010110101100000111110110100101110100110100001010111000101010000110010100000101011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2587[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2587, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100110101101110010001011000010100010110101111100101010100011101101111111010101110110000000011010101111110100001100011101011; 
out2588 = 128'b01111110100011101010101100010110011010110001101100101110110011101101000100101000011110111000100110111010000100111101010111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2588[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2588, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110010000010110100010101101101010010101110110100000110110110001100010011010111011001110010001110100101100110011110010011011; 
out2589 = 128'b11100001100011001100010011001000010001111011010101100111101010001011010111010111001011100101010001011111011111011110011011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2589[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2589, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001110000101110111010001000100110011010111001110010100101010101110001011100100111010111011010100111000010110000111001000000; 
out2590 = 128'b10001100001101100101110010100111100010101000010111001011100111000010000110100110001000000111111000100001011111001010000000001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2590[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2590, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010011101011100111001001101010101000010110000011011000000011101001011100101000110011010101101100010101100110001000011111010010; 
out2591 = 128'b10100010110100000101111010011000110010011011001111000010000100100010110111110110011010010110110101010110001010000111000111111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2591[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2591, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010001100011111100110100011001100110101011111100001100011000100110001110111100110111010010100100101100000010100001110001001; 
out2592 = 128'b01010110110001111101010100111000111001100101100000111001110000110001111001011010001100000111010011101000001001000001100000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2592[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2592, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101011011001011100011110101100001010100010101000101001011011011111111100100001010000001001111100110000011000111000000111001; 
out2593 = 128'b01000001001101111011101011110000110110110011100101111101101101010001100100001111011010001101111000011001001010000110011110111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2593[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2593, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000111111000010010011100111011010110011100111000101100110000010101101110000110111101111010010100100011000000101010010100000; 
out2594 = 128'b01100110001001101000111000110110100101111110101011100000011011001010110010000111101000010001100110100000010110101100110100111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2594[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2594, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101001011101110111000100101100000101101011000100000111011001000010011100101100111010000101100001111110010101001100001010001; 
out2595 = 128'b01110101011101001010010011111010001001101111101010001100011100000011001011111110100101100010010011100101011101011000110011100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2595[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2595, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100001101111111101011000100011110111101001100100101101100010101100111110101010111101011011000101110111011100001111010001001100; 
out2596 = 128'b00000110110111000001000000100001001011000110100011101111011101110001100010100100110001001001110111110101011000000000101000000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2596[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2596, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110010001100111110111010100010000011101011111101110100100110100011000010011010000101101010010010111001111011100011100100001; 
out2597 = 128'b00001001000001010011101110101111010111010010100001101010010110100000110001001100010100110010011010000011111101011111011101101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2597[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2597, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010110111101110001100100110011110001001001111011110101100011000001110101110101111011001111111111001011011110011110000101001001; 
out2598 = 128'b01100101100100000010000001100010110110101000111011111101011100110000111000100100101100100101001011011001000010111010100101010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2598[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2598, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101001101101011010011010100011011101011001101000111010110101011000011101111100101100111110101100010101000110101011010011011; 
out2599 = 128'b00101011010111110000100000000000111000100110100111011010010101011000110101100110001100110101010100011110000000011110010111011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2599[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2599, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110010000110101000100000000100001100100100000000000001111010000011011110100000011011100101011100000001101010000000100010111; 
out2600 = 128'b11000101101010000111101101000100010001010101100111000011110110110001111000010011010100110100001000100111001000101101001000101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2600[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2600, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011000010100110100001010100110010010000100000111000001101110010011101100100001000010110110010110011101010100100011111010001; 
out2601 = 128'b01110100001011011110011010100110010100101010100111111100011001011101010100011101101111010110001110100100010101011100110110110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2601[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2601, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101100101001110100011001100101111001100100011111001010111110010010101000101110000011111111100100011010011010000000100001010; 
out2602 = 128'b01011010100110011100011100001000111101001101000101111110111110111100100011000110000000100101110111001010010011000111100101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2602[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2602, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110000001110110111000100001011110101010000110110110010101100000011001011100010111111000111100010111100010111100110000000001; 
out2603 = 128'b10000110011100011010010000101111001000010001111100010010111100000000100100001000111101000011100110111000101010010000110011000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2603[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2603, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011000111100010110000011001101100111111110110100000110110010100011101111100010110010001100010000111101111111010011111000110; 
out2604 = 128'b11110111010100010100101000010111111111100010000111111011001101000010110110001010110111001001000010001000001011011100111000111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2604[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2604, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110100111001100010011000100011111010100001000011111100000110101110101011010101111000100110101000101011110101001110111101110; 
out2605 = 128'b11000001100110111000110001001111011011100001011010000100110010001011011111011111111001110000110111101110000110100010110010010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2605[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2605, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101010100000011111111110010111001100110101000110001111111001100110101001010101101110000101000100001010101111010010010111100000; 
out2606 = 128'b00000010001010100000011111000010011100101111110111100100100001111100000101100011110100110110100110010100001000000001111110101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2606[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2606, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010100010000101101001011010111010100100000010110001000110010101100111000100010101011111111111101110101011001001100111001100; 
out2607 = 128'b11000100000111111111110010011110111111111010100101100011100011000100011000101100101011001101010000110010011011001011111010100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2607[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2607, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000000111000001111000100100100000010100010110101011001110011010000010000011111110001100000111000100101110000001110101011100; 
out2608 = 128'b10000100101001110011000110111001011111000110100110010001010010011100011100100000100111011011100001111110101011101000110011000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2608[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2608, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100110100001110001101001000011111111100011101010011010001111100110100011101010101000111111100001000111000000101000001100110; 
out2609 = 128'b10100010100101100111101111001011001100110000010010010001001101000101000011101001110011001000101000010101000000110111011011100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2609[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2609, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011001101101001001101111110100001011110100101001011000110010110110000111111010001100010111101010000000011110010100001100011110; 
out2610 = 128'b10001010100111011010101000100000010110011110111101100000100011001110101101110001010001011101110111000100011010110111101010110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2610[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2610, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011111111101101001101011111011000001011101100101000101100100100100111100101011000111101100111111000101000000000000000010000; 
out2611 = 128'b10100001110001100010011010010111010011100000100000100011010000001000011111000110101010011011111001100001110110011000010100111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2611[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2611, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001010110100010000001110110101011111010100101001010111010010100001110010001111010100011100010100001000111010111101011010111; 
out2612 = 128'b00110011010000100010011101010111011111010111111001001110100111000011111011111100010100110000111010010101110101001001000110001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2612[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2612, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110111001011000010000011001110001111100100111101001101011111100001101001100000001000001010100100010001010001100001111011101; 
out2613 = 128'b01000100101110110111011011101011010011100001101011010111011110011111111111010001001111011101101010101100100101011011101111001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2613[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2613, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011111101101001000000010010101000011000100001000100000010110011001010110101010110110000011100101100111100111110010101001011; 
out2614 = 128'b11011000100000001000101101101100000001010101101100101110010011111110100111001110110011100000001111100101101101001101001000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2614[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2614, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111101101101100111000000101011000111110011110100111100101101110011110011011111011001011111001010011101100000010000101100110; 
out2615 = 128'b11000000010010101101001100101100111111111110101000100000110011010110111100011011100000100001010000001010101000101100010011101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2615[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2615, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111101000001101111000000000010111010010111000010111011110111000111000001011000101001110111011100001001101101001011110101101100; 
out2616 = 128'b00001111111000001001000111101010011010000010001100110101011001100110001001001000111100001001111111110111101001000010111101101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2616[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2616, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000100110000010110001001011011101111000000010111111101111000111011100001011010101111110001001110101111001001010100010100101; 
out2617 = 128'b10001011111101010110011111100000000110010001100001010111101101111001111011000000100111001111110011001110111110110110110001000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2617[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2617, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110100001010111110000111001100100001001100100001110001100110110100111001010100001000011101100011110010011000110111111101110; 
out2618 = 128'b01111101011000101110000011110101000000001110100000111001010001010111000000011100100001011010100111000111011000100010000000110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2618[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2618, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110001111011110101100111101011100010011011000011111111101001110111111101110010001100111110100101011010100100000101001010100; 
out2619 = 128'b00011011010011010000010100111110111011001101001010000111110101011100001011000000001000001111110110110111010001011001000001111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2619[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2619, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100011111011011111010110000010000000000100100100011110001000111000001110110111111111011100011110011000110001111000010111000; 
out2620 = 128'b00010111110110110010000110010100010111110011100110010010100000010011010010000010101011100001001110100110100111011000111100001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2620[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2620, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000001001111011111110001101010110011001001010000111110110101111010100010101100011010010101111010101100001011110111000000010; 
out2621 = 128'b00100001000100010001111101001110011011011110000101010101101111110010010111101101100000000101001101111111011001000010101111101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2621[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2621, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001111100001101101110010110001111011101010101001010011110100100000000111110100111101101100110011110110101001101001001110100; 
out2622 = 128'b11110001100000000010111011001111100001100110110011111011101100001001001010001000010001111111001101000000100010111100100000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2622[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2622, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101010101010111011010001110100111001010010111000111011001100110101000000100000110110011100111111101000010000101000000011010111; 
out2623 = 128'b11010000100101010011000000100111001010010001111110000111110101111111111100010110001100100101110100011001001010010110111011100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2623[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2623, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000010000000000101101111001000011011101010011110011000000010000000000000110111111110101100110100100110100001110000011001100; 
out2624 = 128'b00111110001110101111110100010111111101110011000101110001100001000000000100001000010101110101001010111011001100011011101000110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2624[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2624, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100000011110000111110100011110011001111010010111001000011100010100001000001011010001001010111110110011100110100100111010001110; 
out2625 = 128'b11010011111101000010000101100110000010111001011001111011110110000100111001110011010010000110010010111010000110101001101011000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2625[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2625, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001101110111001011110101100010011010101001111001111011000101100110100010111010111110011101111111001010101000010010000000011; 
out2626 = 128'b00100111010110001101001111010110110111010110000000000111011010110101110000000111111011101011100000111011000100101011011101000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2626[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2626, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000101100101001010100000100001011101101001011101110110100110010111011011110110011011001100001010111110101011101001010100011; 
out2627 = 128'b11111001110100101110001011000111011001101000000111010001100010111000101110111011110111100010010111111101000001110000110101101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2627[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2627, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100000011111100001001111100110010000110010011000110001011101101110110101001001000011110110000011000100011110111101000011000; 
out2628 = 128'b01001010101111101111101001111111011001010011000011100100101011011101100011010001110000010101001011111110001111001001011110100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2628[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2628, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011010011010111100010100110101000011101000001111110001100001011110011100110011001111111100011111000100010111100100010101001; 
out2629 = 128'b01110101111000010111011100001011011000000101010110011001110111010010111100011100111100110000100101000010110110010010101001010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2629[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2629, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010000001110110100000100001010111111010010111111100001101110000110111011100110100001011110011111110001101101010111011010000; 
out2630 = 128'b00000100001110110010011110010000111111001111010101101001101010010001100010011011011000001111110101110010011101010010001011000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2630[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2630, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100000111101010111011010101001000111010011110101001010001110011010111011111011010010101100011000111100010010111100011111110; 
out2631 = 128'b11111001011110011000000000001001101101001001111010010010010101101111000000100010001101000111011011111000110001110011110100101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2631[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2631, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001101100100010100111011110000011000100010101101011011010000010110101000010101000001111001110100000011110100110100100101001; 
out2632 = 128'b11100111100101110111001010010001010111101010100011111111101110001011011100010101011100000111011000100011101010100010100011010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2632[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2632, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100000110111111000000100001101111010010011110100011111001000101000011101101010100110010000000101101110101110100111110100010000; 
out2633 = 128'b11110111001010110001110101100101111111100101110110000101101011010010110011011010110001111101010011010011010001100001110100011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2633[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2633, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111000010001101010111001001000111101001110000010001101100101101111111011001100111010101101000011110111010101000011111111111010; 
out2634 = 128'b11001001010001111100001101110100000000101111110110101001111111101100000001111111101111110101010001111010101000101011010001100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2634[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2634, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011011111110110010001101000010001000101000010110100111100010101110101110010000000100110010101011110010010110100001100011100; 
out2635 = 128'b00011111101110111100011001100111010110100101000111011111100000010100011101011110110010000111101100000010001000110110010001100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2635[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2635, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001011101001111001110011101111010101000101110001010101011000100011100101111100110011011011100011111100100100110111010010100; 
out2636 = 128'b11011000011110011000010101010101110101000010010011001010100001100001000011111100111101000011101011001110111100000010101101001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2636[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2636, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101010010010110000001111011110000000111111010010010101000011100110101111010010100100001100110001101110010000101001001010010; 
out2637 = 128'b10110001100001010111100001101111101110001100000111100011001010001000110011111001100101001000001100100000011001101011111000001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2637[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2637, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100000111011110111110101001010110110101001001000001111001110001001101011011101011001111111010111001101100100000010010010001; 
out2638 = 128'b11011001011001000100010011101110110111101100111011100100100001101010100000100001000011010101111011111101101010101101111010100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2638[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2638, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100100001011000010101100111101111011000101010101110111110111110011111101111010000011111011001100101110000001100000101011111; 
out2639 = 128'b10100011110011101000100010110001001010001011111111111111010101111011011110010111110111010111100000000001110000100110110010001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2639[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2639, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001100010100010011101101010011101100111111100010111010010100011001110101111110011111111101001011111101111010001110010000100; 
out2640 = 128'b01110001100100100000010011110110101111110101011101011010110111010101001010110001100111000101000000100010010011001101110001001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2640[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2640, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011101101010000110000110101010001100101000000011100010000111000011100000110000001111111001010011001011100001000101000110000; 
out2641 = 128'b01011001010001100110000010110110110001100000001110000100010101111111010011101010100011000000110001110110000101111000010100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2641[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2641, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101010000001101010110101011000111101101001110111100000001000001001100010100000000100001000110100100110000100011110111010110; 
out2642 = 128'b10000111110000111000010011100111001001011010100010010110001001110000010101010001000100000011100010001110010101010111010110000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2642[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2642, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010100000111010011100000010111110010110011000110100110110101001100101111101011001100011100010000110011000000001111010001011; 
out2643 = 128'b11111101000100110001110010101111110101110001110101001111001011001110010101001010000111011110100000011101011000101101101001001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2643[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2643, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010000100100110010100101001011010011000101001100100011001111100101111001001100101011000101111000001111001001010100101001000; 
out2644 = 128'b00110001000101001000110101100011000001010001110000100000110010001000001001111100011010011100101010010011101101101100000101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2644[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2644, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101110100001000001010111001100010010000011010100000111010100100011100110001111011100101100001101001100110001001110001100110; 
out2645 = 128'b11100111100101010100000001101011001100100110011011001100001110011101101000000111001100100000001011000111101010001101011101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2645[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2645, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101000001000100010110110110110011011100010111011010000111110111011001001101011110000001010111100011010110011100111010100001; 
out2646 = 128'b10101100010110111001101010111010100111011101001001010001100110101000000001001101100001110010110000101110100011110001000011101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2646[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2646, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001000011110000011110010000111101011100110010111010110000001001011100110000111101100010010110101011100011010010111111101000; 
out2647 = 128'b10011011100101100101101101010011000010101111110001110100110010111101000100010101010100110001010000011000100110100011100010000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2647[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2647, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100111011011100001001010111111001000001000110110001100101110101111101110101101111100111101111101001100001101111001100000100; 
out2648 = 128'b01010111011001110101011011110111111100101000011011110110110001011101010101000100001011010011110000101101111010110010001100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2648[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2648, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010011010000100011011101111000010011110000010011111011011101100111011101001011111000100000010001111110111100011100001111010; 
out2649 = 128'b11010001000111111110110010100100111010000101010001011010010111011011011011101011110011110010000110100000110011000011001111000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2649[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2649, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000100010001111101001110010000011111100100110010010011110111011100011001111000110000001001101110010110111100000110111110000; 
out2650 = 128'b00101001001110011100110001011111010110011000101111110001111101000010010000011111001010001110001011000100110111110011000111101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2650[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2650, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101111100001001101010101010100100101110100010110001010101001100001010110100110001010010011011101000100000010110001110111100; 
out2651 = 128'b10110000110111110010001000110000000110001110010010000001101011110000101111100000100001011101111111010101101010001000011000000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2651[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2651, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000011011110001010000110111111110011010001110110001001001011001010110100001011110100010001001001101000110001101011110000110; 
out2652 = 128'b11110010110000010001010100000100110100100111010011010110100011001101111000101001000111001101100100111010010110100000010001111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2652[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2652, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010000001100000101001011100010001100110111010000100011011010001100001001111000001101001010000000111100001101110011011110001; 
out2653 = 128'b11100001011000001111010001100101011010010101011001110010001101011010100010110011001001011101011011011100111000111100001000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2653[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2653, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101000010110100000011010101011100000000010000011000101001000011010001101011100101011000100000101101010010101000100000010000; 
out2654 = 128'b10001101110101001101001100001010110001010111010110111001001100101011111000111000111010011011001111101010110111000011000100001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2654[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2654, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110000000101000000101101001100010010011100110000101110101100001011101110110011010101111001100011000010111100011110010000110; 
out2655 = 128'b01001101000010110010011100110000110110101101011100110010011100000111001010110110100001101100011010000000011110000010010101001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2655[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2655, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101101011111010011000100011010010111111010111001001011010110100101001001011000110011011100011111010011001001001011001010011; 
out2656 = 128'b10000100101101011011011011111111001100100111000110101101000010011111101110010101000111001110111101010000001101011000000011011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2656[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2656, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101010101111100000101000010100000101010100001111111000001100101110001111011000011101010000001011010101110100000101001111111; 
out2657 = 128'b10111111100111001110001101100010000111010111000001110010111110010000000001111011110110001101101000100011111001000100100110100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2657[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2657, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001101110010110001011011100000000100111011000101101011010100011101010011110010011111000010011110110011000111011001100101100; 
out2658 = 128'b10010000111100100001000001000001010000100111011101100101011000111111110111101010111101000100011000101110001010111001011110011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2658[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2658, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001010001000011001101111010011111011001001011100010111001000101111001110010001000001000000000100000011001010010111110011100; 
out2659 = 128'b10010101010100000001110100010110011110011111000000000000100000101110000010100011101111001000101010000100001111011010011001100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2659[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2659, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001001001010111110110011001000111001110011011100100111000011000110100001101000011100010010010001011100111010000011110011010; 
out2660 = 128'b11110101010011111000111001111111000010100110001000100111101000100101100101100111000101000110011110111001110100111111110000111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2660[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2660, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111011010011010011110110001011101111100001100101001010100000100111110010001101011100010011000011010000110111101001001001001; 
out2661 = 128'b11010011100011010001001110101000001111101010101001111100011000011010001101101110100010010100101000111100001111011110000011010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2661[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2661, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010101011111100001110000001110110001010111100101000110010000010000110000000010010100011011110101111011000000111001101011111; 
out2662 = 128'b01001011001011011101000110011100001100000011011001001011101111100001110101110010000111011010001001100101001011011101110100111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2662[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2662, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011100110010010111000001111100100000100011111010000110100011011000111010101010011011000001010011111100100100011100001011001001; 
out2663 = 128'b00101011111001000100100010111101011110100001110101100000111111011011000100010110110010001110101111001011001001010001111001011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2663[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2663, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010110010001010010011000111110011100011100110001100001000100010010000000010110110111111010000110001010100001111011100010110000; 
out2664 = 128'b00111100000011111001000101111100101100100000100000010000001111110000010101110111100111110010010111111001111011001010111000000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2664[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2664, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101101001010010010001111001001000101100100011111110111110100010110101010010111010011111011001001001001111010011111101010010; 
out2665 = 128'b00100111001111110110000000011011001100000101110101001110101100011101001111010110011101110001001111110111101111111111001010010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2665[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2665, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010101101110001111100111010111111110001011001010100111011101111011001100000011110010001001011110010101010111111110110000011; 
out2666 = 128'b01100001011001001011000110000011111010111010110110100100001011101100111110000101011011011000101111001100001100011101000101101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2666[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2666, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001110101100010010101011000111010010000110010010110101111011001111101010001100100100100010100000011110100011010110110001111; 
out2667 = 128'b11000010101011000100010011110101100001111010000110001100010001111111100001011100000111000111111110101100110111111100111111001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2667[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2667, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111110100101111011000001011011110111001010110100100111000010010111001101111111101110001101111010100001111111010110100111110; 
out2668 = 128'b00100000110010110111011111010010011100110011110110110001010000011001001111001000101101100011110011101001101010110011100100011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2668[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2668, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100110111110101010110001100010111110000111010110010010010000111001110110001001001011111001101101101101101000011111011011011; 
out2669 = 128'b10110110110101011110110110111100101110001000011110000011010010001001110010111110010010101001000111100011001100001001110011100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2669[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2669, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010101000000001000101100011010111011001100001000110110110110101000001101010110010101100101111001010000100000100111110110100; 
out2670 = 128'b00101101111101100000010000111111110010100010111111101011101010100010001111111010011101001111110001110010110110101010010101001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2670[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2670, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101000001101110111010100111110111110011011010111111101101111110100001000011000001110000111001110111011100000011100000100111; 
out2671 = 128'b10100010000010101010000111011011001101000000010101010111100010001001101101111111001111011000010010101000110101111100101110111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2671[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2671, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110001011000111011011010100010110010011110010100000110001011011110100010110111110101111101011001000101001010100001011101011; 
out2672 = 128'b01101101011100001001100101100010011101000011110100101110011110110001011101111111010101001000000010010101101111111110100111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2672[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2672, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100000000110001000000000011100011011111110110011001111001101111111111000010000101100111101010001100001110100011000110101110; 
out2673 = 128'b00111110111110110000111001100010011001110011100010001000111011110000101011110101010111000101010101110101001111110010011110010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2673[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2673, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110011100001100110110100111011000000001100010111111111001000101110010111001100001011101110001100011111111011000110001000011; 
out2674 = 128'b10101010101110011010001001100010110110000011000001011101100100110011100001110010100100010000010011100110000000001110010111101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2674[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2674, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110010110111010011000111100001010010000100010111100000001000010001111100111100100010010101010111001111110001100000011101110; 
out2675 = 128'b11001011101010011001001010000000000010001010111001110011111101110111010111110100010101001011101010011110001111101111001100111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2675[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2675, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101110011100100010001111010000100111101110001001100001111111101010101011100001001010000111100010111101110111110010011000001; 
out2676 = 128'b00001111101010011110011011110111111011001100010011111101001010000000011010111100110101101011000000101101000001001001100110011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2676[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2676, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010111011111010000111001110101001110111010000111100100001110001000000101101110111100000101111010101101111010110100010100101; 
out2677 = 128'b00101001001101000101011000001111010000001001000111101001110000001111011110110011111110000110001111011011001011101001001111011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2677[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2677, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111110111111000110110011000100110101111011000101111100100111110010110011111110001011100111111111111001000011011101011110110011; 
out2678 = 128'b01011101111100000010011111111110110110011110011110111111101110000011111100010000000000010011001101001100001000011000111000011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2678[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2678, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100111011011011100001100111100110011010110001110010111011000001100010100111010100010011000000111110110110101111011111100110; 
out2679 = 128'b01100011100100001101101001110001110100000010111111011101100100110101110100100011110001101111010010010000000011110010110001100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2679[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2679, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100001111010110010101100110010100101010001010101011011100100101001101001110011100111001011010100101011001011100011100001110; 
out2680 = 128'b10001101000110110101000101000001011011101101110000000111011011110011111011100111011001001100011000010111000101101101100000110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2680[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2680, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110010111010100110011011110000100010001010110011010111100001001000111100000110010110001110101111011100100001011001111011000; 
out2681 = 128'b00011110010001010000100010010000001010111101111000010100100000000101001101110110000010101101110001010001010001111101000001100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2681[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2681, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111101100101010110111100110111111110011001011011111100001110101000111111100010111010110110110011100110000000010010000010111; 
out2682 = 128'b10101000111001001100001011000101000010000101111110000101101010010110111110110001011001000100101010011001101000010101111110100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2682[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2682, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011110000100010000100001111011000101110110101110111011010011000000001000010111100100011011000011001110111000011110110101001; 
out2683 = 128'b01100101111100100000010101101110100011110100010111111111011011100111100010101001100110111001000011101011000111100101010110111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2683[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2683, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101100001100000010111010110001001100100111110010111111110000100100111000000101101110110100111101111001100111000001000111001; 
out2684 = 128'b00100110000001101110000100111011010100100010010001101001000101101100100010100100101100110100100111001001110101110011100010011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2684[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2684, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001010011000101010101100101100010101001111010101001100100100000010110100110001001011001101110010111111101100101010001111001010; 
out2685 = 128'b11011001001000000110010100111101010111110110001011011011111101000110011101001000000010110010110000001101100010000010001010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2685[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2685, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100000110110011001001011000000111001100101010000101110110100111110000011001100011010110001100111110110100101011100001011000; 
out2686 = 128'b00100111111110110001110000001000110111011111100000110101000001000100101111010001010100111001000110000100101011100110101000011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2686[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2686, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111110001000101000100001001111000100000010010111100010001100011011111111100010000100001101100111100000001101000100000011001; 
out2687 = 128'b01101001111010111000000010111100110001010110011000001100101101100101100110111010000101110000000010100001110111011010001010010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2687[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2687, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001111101110001000110000000010010101110000110011011101111100010110011000111110111110100101111011100110111101110001110111011; 
out2688 = 128'b11100001010001000011000001111110010100110100100110000101000100100101011110111001000100010000110010001101101010101100010001011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2688[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2688, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100100101010111111011001100111001000101100111010110110100101111010000001001001001100001110011100001110000101110101001000011; 
out2689 = 128'b00010101001101100101111101101001010110000010100100000000111000101101011101000111100111011010111010011110001001011101100101001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2689[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2689, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111000110101001001100000111011101001001000000101011100010011110111100100000100011010011011011001000110111001010000011110010; 
out2690 = 128'b00100100010101010100101011000000001110101001000000101101110101100010110011101011011001110110111010101100100111000011110110110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2690[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2690, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001100000110111101110111000100010100111100100011111101001001110111000100111111100100110110000000000000111101010010100110111; 
out2691 = 128'b00110111111001101110100011001101010001011111110101011011011001001001000011000110010110000110100001000010101011111010010000100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2691[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2691, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110000100110101010101110010010100010111110000001100100110100101001010011011101010000001101000010101001100011111110000110001010; 
out2692 = 128'b10110100000111100101101000111000001100110011101110011101111001010010000011000110000100110101000011001110111111111101111010001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2692[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2692, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011001001001100101011000010101100100101111111111011010111001101111000110000110010111011010100001000100001110110000001001100100; 
out2693 = 128'b11101010000000010101110010101011011111000000000110100100110000000011010111011001000010010101010011101011010111001101110010010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2693[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2693, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101001010111011011001010011110010101111110011001010111000100010101001101101111111100000001000111001110001011101001101110101; 
out2694 = 128'b11111100001011100110110010001000101010010100001000111110110010111001100110111111110001100110111110110101001010101011110000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2694[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2694, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111001001110010011010101011111101111010000111111111000010111010000101111110010000010001010010101010111010011000101100010011; 
out2695 = 128'b11011000011100101010101110111100101011000111110111010101010001000101110100011100010100010111110110111100110010100101000111001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2695[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2695, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111101111100010101001000001010000111111111111110100010100101101000101010010110000100101010001110100011000011001110101010011100; 
out2696 = 128'b10101010001000010100011011101110010101011101000101111011101110110001010001100001001111110001011101110000011110100111111010011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2696[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2696, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001100001101010101110111000001110010111001110001110001110100111000011011000100100111110111110100100101110000001010101010010; 
out2697 = 128'b01010101100010011000110100101011010101001010111011011011000100011110111111011000111000011101101101000011001100110000111111101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2697[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2697, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111000000100101101101101000111001011110010101000010101000110100111110110101100011001111010010011110001101000100110010011101; 
out2698 = 128'b10011001110101101010101010110000101101010101011011110101111010100010101011000000001111100110011000001100011001011101110111110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2698[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2698, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001110001011001010110100100001000010101110001010001001111111011100100011110001100001001101000001000011101001100000101110001; 
out2699 = 128'b10000010100000100101101010010101110000011111010000011111111101000111101110001001101101100000110111100111100011101010000101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2699[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2699, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100110001000100001001001010011001000011001000101011001001000110010010100000010000010001001000001111100110000010110101101000; 
out2700 = 128'b10001001110001100011011101010010010101010100110101000011101100010010000111111011110000000000010110010011100111110011111011101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2700[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2700, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100011101000111111100111100100100000011011001011010011100000101101111100110011011010010110011011110100001110111000011011110; 
out2701 = 128'b10001011010001101001001001001000011010000100001010101001011011110011100110101000011110000001001111000010110000101111010101100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2701[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2701, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111000001100001111110010000100001011101100011011000101110110001011101111100111101110010110000110001101100101101011111100110010; 
out2702 = 128'b10100110110001010000101100010010010010110010011100001100011110101001101000001001101110011101110110101110011100011000001110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2702[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2702, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110000101001100111000110001100011001111010000011011000100100000011010110111110011010110110001000110001100000010100011101110100; 
out2703 = 128'b00100110101011100011111011111010100101001111100000100110101001111001111001001010001011101101110001110001110111000110111001110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2703[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2703, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111111100111110111101011100110010001011001001110011100100111010001010000111010111101111011000011010101010011000010111000101; 
out2704 = 128'b00001000110110110011011101000000101100111101010101100110000101000110110110101000011010000110000010111011100001110100110110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2704[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2704, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101000010111111110001011011110000001101001011001100000000101010110000010001100011111101111111010111101000110010101010100110; 
out2705 = 128'b11010010001101010110000100100110010011101111010001100111111000111110011000011001011001101110001101011010101101011001001111010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2705[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2705, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110000000100111100000011100100100011010010100011010101000100000011000001000000010000111101001001101011100101111111011011101; 
out2706 = 128'b11011001011000010110111100011010100010111100110100101110010110110001100010001011101111111110011101011001110000100110000000110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2706[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2706, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111000110001100110111001000001101101011110010001010100101111100110000011101111001100101011101001001100010110101111101001111; 
out2707 = 128'b01110000110100111000110001001001010110010111000010100110000000011011101000011011100001001010011101101111110011010110010010111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2707[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2707, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001000000110010010001000011110001010111000101111110100011011100110111011100010000111111001100011111110100010110000000001101; 
out2708 = 128'b00010111010010100101000000000111011011000011101000101110010101011001111010110010111000011001100001110100101100110010110110010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2708[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2708, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111000101111001011111011111000001000001001101001001111000110001010011111010010000111101010110011101110110110110110001011011; 
out2709 = 128'b11100100000010101010000010011000111101000010001100001000110100111111010110000000010101100110111110111110101110011100111011111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2709[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2709, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000010111110101010001100001110011101000001101111000101001010011011100000100011000000110001001000101011001011110111001010100; 
out2710 = 128'b00000100010001100111011100100101111001010010000000101100000001001110110001101011111001110001000010110110100011100001111001111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2710[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2710, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011101110111001101001110111100011010000111101111100100110100111001010110001110010110100011111001000111000000111000110110101; 
out2711 = 128'b01100100111100000000110111101011010010101101001011010011010010101011011010111000110101000100101010111111100110111001111110011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2711[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2711, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111000001011111110101111000001010111000110111001110110001010100001100110010100111110011110100110111001011101001100100011110; 
out2712 = 128'b00100100001011010111100101110010010011111000100011001000011101110011110110110111011000111100000110001001110110111101001000110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2712[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2712, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011111101000001101111011100001110001010001100101101110101010010100000000001101001101000110001001111010100000111110101011110; 
out2713 = 128'b00101001110101101011110010101001111001110110101111001111111010001111111101010000010001101000011010011010011101000111111100111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2713[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2713, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011011100011001011100101001010110000000101100010000101110011000110100000010001000011000101100110010000101101101010111011110; 
out2714 = 128'b10101000000100000010010100111111101011010110000111111111110101100010111001100110100100100000010010000111011011001001111011101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2714[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2714, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000011111010000001101110100110010000011001100111110010110011111100111011100100101100110011001100010010010101001011001010100; 
out2715 = 128'b10001100100000000110110011110001101011001101010001011011011000011111001110111011000010101001000001000111011111010000100111110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2715[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2715, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011010100011001101010000101111011111100101101000101010011100000110000110110001100110011000100010001010100001001001100101100; 
out2716 = 128'b00010001011011010000101000001110010100111011110001011110100111111111001000000010001010100101000100101010010110011010011011111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2716[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2716, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110010011011000010000100100110110101111000011111011110010010100011110011001001000101110110111101110000111011110100011110101; 
out2717 = 128'b10001000011000101000111101100001110101001110000110000011000100100110111001101001101110000001011100110100001001011101100111011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2717[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2717, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100111111010011001111010101000101110000000011110100011010000100011000111011111010011101001000000101010000000111000011010110; 
out2718 = 128'b00100100100111100110010101011000000011011111000011001011010000101000100010100111110101010010101011010100000101111111110101101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2718[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2718, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010011000000011010101110100010110101111100010010010101001010101011001101000000111010011001010011101100001101111100100100011; 
out2719 = 128'b00000011000100010110000000000101010111011101111111111010110110101000010011000111010010000000101111100101110001011010110101000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2719[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2719, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110010110110010110101111100100101000001000011001101111011101101101001110100101111000101010100101111001110000111100101010001; 
out2720 = 128'b11000011001011101101000110110001100101101001110000110011100011001110101010011001010000011101011101110100010011011001001101001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2720[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2720, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000111111001111101001011000101001011100101111001011010011000110010011011001100011011010100010000100110011101011000100101110; 
out2721 = 128'b00100000001111100000101001110101101000001010100111000000111011001011111001110001111011010011011010001011000111010101000110100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2721[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2721, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101010100101100001111010010111000100111111010100111111101111011010101010010011101010100001001010001010001000100001011100010; 
out2722 = 128'b00111100000010101111011101101000111010111111010111010111000101000101110011010011100000111011101000001010001001011011001000000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2722[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2722, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011101011000011000111101010101100011100101111001100001000101010110010001011100100011101111011110001111010000111110011101011; 
out2723 = 128'b11010100000110101010101000001001110000000010111101010000100001111110000110110001100110000011000100010110100001011101110000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2723[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2723, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001111000011101010100110010001010010110101101000010110100100001010101011110000100101100110011101011000111100110000001010101101; 
out2724 = 128'b11001100011111010100010111011110101010110011001011101100001101000000100001111110011011011101001010001101100110111011001010001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2724[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2724, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110100111001110101001101010010011000111001010110000010110010001001010111100001101001011100010111010100000111000010101011110; 
out2725 = 128'b11110111010010011000111111000100000100000100100110110101111100011001101100101110000010101000011001110101010010100001110100001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2725[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2725, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100011010001000011000110110110100010011001000010111010011111101101111011110010000011101101100011100001000111010100011111001010; 
out2726 = 128'b00100010100010000101011110111100111110001100100111110011101111000110111001111110001010110000000100111100111001101010010100000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2726[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2726, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011000010010001111111010000110101010101110110100101011111110001000010111010001110010101100110011011001100111100010111111011; 
out2727 = 128'b11110100001000110101101111011101000101101110010001101111101000010111100011001100101001000101111100011100000111011010110010101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2727[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2727, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100110110101110111100011101111111110101110101000001101101001011101111010010001111110000000111110000100100100101010001011001; 
out2728 = 128'b10100000111011111011011001010100111110011011111001110101010100000010100110100010011110100011101101110000000011100100000110101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2728[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2728, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111000001011100000010000000000010001110001000010011100110101111001000101010110111011111110000000000011001100100000100000111; 
out2729 = 128'b00110100011101110111000110101101010101011111000100010000111001111001000011010011101110111000011011001010100101001001000100001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2729[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2729, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010111000110000010110011000110100100001111001001001001010011101010111011110001000000010001100010110111011011010110110011001; 
out2730 = 128'b11100011111001010011100010110110010000110011001110010001000001001011001101010000001000000101111010010011000011100000011110000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2730[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2730, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000110011011111101001000101101000000100110111011101101001000111000110101100011001111001110011000011001001011111101001011111; 
out2731 = 128'b11110001001000010011001001111001001001111001001110000010110110001100010101101101100101111111111100110001101111100110000101001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2731[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2731, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001100011011100011010000010001101100100110001011110001011010010101101000001011101010111101011010011100000001110111000000010101; 
out2732 = 128'b00011101101010011000000101101010001101100101110000010111000101011010001110101110011001001110110111010111101100010011100110011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2732[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2732, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101000111001100000111011001101101110011000010110110111010010000001011001110010000011000110011000111001101010011100100000000; 
out2733 = 128'b11101011110001010010101001111010010000001010101111100000010111001111111110111000000000101100001011010011111011010010001100101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2733[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2733, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100010001010001100000110100010111110111010011000100100001111111011100111010001010100000010101101111000111100111001100000101; 
out2734 = 128'b10001011110000010000100000010001101110101011010100000010100101000111101011010101010001100010010110110010101100111110011001001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2734[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2734, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111100010001001010101101100011010001000101110110110111000101011111100110011111010101111111001101011001101111000000110010100; 
out2735 = 128'b10010111011110000110111000111101000010010110010111010010011000011110010110110001011011100100111000011111101101100101111000110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2735[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2735, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111000111110100100001100000010000011010010111101101011000100001010111101011110111001111001110001111000011011010011111000001; 
out2736 = 128'b11100001100010001001011000000100000111110000100100111011010011111111010001011001111111100010100111011101110111011000101011111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2736[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2736, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111010111100110010000011111110001111000111010101001100100101001110111011101000000011110111011101000001100010011111100100101; 
out2737 = 128'b11011100110011101110100110110001110111110101101101011001000111010100101101000111001100111010111000010010111011101100111110110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2737[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2737, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000011001010110100101100101110110110010101011010111001101001110111101011000101110111001001010001100011000110001011011001000; 
out2738 = 128'b01111010110001101111101101100111000000101000010011010110101110010010110001101101010111110111011100100100001110000100101100100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2738[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2738, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100011100100101000101110011111011100001011100100101011101111101100111101000101010101111011000001111100010001000010001000010011; 
out2739 = 128'b00110110000101100101110100110011000001011100101110101110011010110011100010011010000010111100000110000011010111110001010111110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2739[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2739, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111110100000001001000100000001100110110000000101000100001011001010111101001001101101111110111011010111111111000010011101000; 
out2740 = 128'b01101100100001101100000101001100011110101111111100110011001011101101100001101000100101111101111101101000010001101000101010101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2740[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2740, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010101111001110001001011111110101001010110010101011001011111110111100001100001101000101010000001110000010101110110000000001; 
out2741 = 128'b00001111010101010010101001101011110011010001100101011011110111000010001000110100011001001111111101010111101001101010101111001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2741[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2741, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010101001110100111010011100111001111100111010101100000010010000110011111000110100101011000110000000010111011011010100100110; 
out2742 = 128'b11000110011011011010001111010110011100001000111000000111111110101001000010011001111001111111110001011011001000111111111001001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2742[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2742, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000100111010010010001111101111110101000010101010111000100011110101001000101100101001110110011001100111101110011110011010111; 
out2743 = 128'b00010101010110101001110111110011101110111100011110001000001000110110110011100101001110011100101100101001000000111100100001011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2743[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2743, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000110010000000001111101001000001111111110100100011000011101101000000001100101010101000110101101000111101000101111111100000; 
out2744 = 128'b11100110110000001110111111111011110001101011101100101011101101100010011011100110101010111110100010010111011010111001111000110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2744[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2744, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111011010111110100110101001010111100010001101111010101110111010110111110101000000011011001010100000110110000011100000010011; 
out2745 = 128'b00011100000111110101101110100000110011010011011100100110110001011001111100010101010010110001010011000011101011001100100110001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2745[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2745, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011111011111001111100001111101011111101010101100000010110111010011010110011001000100110111010001111100111100100010011011011; 
out2746 = 128'b01010010010000100100111110111101100011110101111111011100111000110001000001011111101111011110110000000010000110001100010111001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2746[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2746, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001110111111011101100001010010110011110000100100011000101001101101110110000000101010010100001110111100011101001000100001011; 
out2747 = 128'b01011010010111111011110001101001000011011111111110001000110001110011111100111110010010110011001100001100000110110001111111010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2747[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2747, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000001010100110001001101001111110011100011000010111000011111110110001011010000110101011101001110011010000101010100101101011; 
out2748 = 128'b10000001100001011110100000110110110111111010011000101011100010110111101111111000100011110110100001010001001111001101101000110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2748[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2748, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101111110010111100001111100110100001111000111010101000111100110001101010110000011010011000010100101101000001000010001110111; 
out2749 = 128'b00001110001000011110010000100001000110001101001110000001001011011001010100000000000111100001111111011100011001011000110000001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2749[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2749, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111111010011001100110000001010001101100111101011101110100110100110000001110010011101000100101000101110001001100011111100011; 
out2750 = 128'b10011110101100010110010111000111111011010111111000011000001011000010110001101111110100001100010011010100011011010110100110011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2750[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2750, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110101101001110110100011000000000000100100001100110001100001110110000001001001100110000010100101000101101100100111010101111; 
out2751 = 128'b11111110010000101000011000011011010011110100000111010100111000001110111110010010111111000010111111010101000110110111110011011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2751[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2751, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010110111011100110000001010101010100100011110011111001110111011110010001100001010101100011011100011011001100100001110110010; 
out2752 = 128'b11110010001001111100110100011000010011100011111011011010011110001111010010010110011000001001011101001000011001110110110101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2752[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2752, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011110101111111111100001000011100011110101011011001101101101110110011110000000010011010000100000101110110011110101110101111; 
out2753 = 128'b01010000000000101100101110000010011100111000001001101100111010100010100101100101100100100100011110110101100010111111101010100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2753[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2753, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000011100101000011111101111100111101101000110101000010110111010100100001011000011000100100010011011010111001001101101110011011; 
out2754 = 128'b01001000011101111000010000001011011111000111100101000110101010100111100100100110000001001101011011011011010000000110101100111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2754[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2754, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011001101010001111100111101011010110000110111010001000011000010010010101110111100010111010111100000011111110011100010001101; 
out2755 = 128'b01110010010100111111100011011111010000110110100110011000000010101011010011111010100010111001010101011011101101000010000001001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2755[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2755, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011000001000100000011000110010001111110111011100110110110111000100101000111001010011000011001101001010001100000011100001000; 
out2756 = 128'b11110111110000011000100011000000111111011101111111011001110001110011000110100010000110011011001001011000101111011111101000011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2756[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2756, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100001101000010001111001110000110110000111010110111011110110101100001000000011000011100111001001000010110110010001001001110; 
out2757 = 128'b00011110001010000000100000001011011101000011011000111010010111101000010110111110110011110001010111101110111110001011110100101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2757[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2757, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110110100001101111110111000011000001111110010001001010100010001000000011100001100101000101011111011100001111001101111111110; 
out2758 = 128'b11011100001100101010111110010000110100101110111110010111011011011011100111100011000000000010011100011110000100100111010101011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2758[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2758, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010001011100110111010101101111110110100111011110111100011000100101001001111000100001111011110000100000101111010111111111101; 
out2759 = 128'b00111000111001111111111001011111101011111001010011000010011001001110010010111010100110100101001101011001011010011000110011100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2759[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2759, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110010000001011010101000011011100001010010000011001001010111100010110011011001110111111111010000110100001101001000111000011; 
out2760 = 128'b01110011011110011101111011110101111100101110001001001100110011010011100001111110100011011010010001100100001011101101110111111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2760[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2760, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001101100101001011001000011010110010111010011001100011101110110010011001000000100111111101101110010010001001000010101110010; 
out2761 = 128'b01111110110101100010011010110110101110111000001010000000100100011100010111101001001000001001001001001110000111110001100010110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2761[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2761, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010010010111000010011000101110000010011011101111100111010010000011101100001011111100011001100100000011111010101001010010010; 
out2762 = 128'b00100010011110110001110100010111110000000011111010010111011010100010110101100100111011010000111011101010011001001010010001000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2762[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2762, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110111011011101010001101111011101101100011010011101001111110101111000011001111101011001110011010000011111100111110010010000; 
out2763 = 128'b10011011000101011001101001010110100110100100111110011111011000001001101010000010011010110001011100010011111110010111011111101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2763[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2763, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100111000100010001110010101001101011011000001000010101111010101111111001111010010110111100000010101000000110101110010111111; 
out2764 = 128'b10001001111001100000110111000000110101110111110011011100101111011000101101111011001001010001011011101111111111100111001011100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2764[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2764, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000001001100010100000010101111000100100110111111001000011000011110100101001101010111111101100011101000001001100101111101110; 
out2765 = 128'b11100011010011100010000101110111010011000011110011100010100001001101110101010101000011101011111101101010100001110110010101011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2765[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2765, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111000110111010101100110010100111110100001001111101110000011010010010100000001000011001010001111010001100000011111010010111; 
out2766 = 128'b11010101101001011111110001101011001010110010111110110001101111010101100001000110000100001010001011101000101110011011111110000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2766[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2766, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011111111001101110001001110000100000001000101111100100010011000001010000111001100001111100000000101111000001101110110101000100; 
out2767 = 128'b11000000100110101101010100110001110001100100000001101100100101000111010010010000110010100110001111011111001001111000000110100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2767[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2767, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001000000101101111101101111110000100001010101111010100101101101001001000111100111100000000011110011101000000100010001011010011; 
out2768 = 128'b00011100111001101111110100010000011110100111001000000001010100101100001101111011000001010011110000010001011100000101101100000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2768[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2768, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011010110111010101100011110101101111101001010001101111110100110011000011111011011111010100010101001101001101011111011110000; 
out2769 = 128'b10010101111000000101010001000011111011100111010001011101100100011011111000010001010001000101001111011110100111111011100011011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2769[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2769, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010010110010000111010010011100011111000001011110110100101010011101111011100101100110100011111010011001101010111111101011001; 
out2770 = 128'b00110111101010000010010110110100111110110000111101010000101000111110100001011111101001010101011011110010010110100010100010100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2770[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2770, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100000111001111000101100101000000111011111000100000101111110001101100011011000010000110101100111110111110001111010001011110; 
out2771 = 128'b11110111100100101100001000011100110001010011010100111110001011111010100000111011011011111101001011010111101001010110001011100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2771[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2771, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110110001111001111111011001110000001000010101110100011001100101111111111010000001100001110001010001011000101000010100001001; 
out2772 = 128'b01110000101110011000001111000100010101110111100011000100101101001001001000010011000001100010011010011101111100011001100101100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2772[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2772, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111010001100001100101010000001111000000011101001101000000110111010000010001110100110001010110101001111101001101000101010100; 
out2773 = 128'b10100101011110011110010101101010001000011010110110010111011000000100010110011000110001111101100101100010011101010110101000101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2773[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2773, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100000000011010011001010010000100000000110000011011000110001111101101010111000110100010001110001000011011101111001000001100; 
out2774 = 128'b10011010100111111110001011000101011110100111110111101010010010000101110111010110011001011100101011010111110000010110001011011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2774[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2774, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011100100000000000001010100101011001101000111011101000001110101000011000110100100100001010011001100111110101000001101111111; 
out2775 = 128'b01111110011011010001011101100001101000100010000001000011000110010001001001000001110011010011110000110011010010001010011010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2775[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2775, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010110110101110110001011000000110010100101100011010000100011000101101111110101110010011011111011111010101100011111000100001; 
out2776 = 128'b10100000001110010011111110000010011111000101111110010110100101000100010010111010001100110011110000001001101001010100110010011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2776[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2776, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010010100101001111110111100001101000000100100010111101000110100011101100000010110101011100011011000011101100010000100101111; 
out2777 = 128'b01000110011001001110101011001100001101100110001001110101100000000011100111101000111111001011111110101010110101110100011011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2777[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2777, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000010110011100010110001011100111000000001101111001011100001101000001000000000010000000101011010001010111101010101111000111; 
out2778 = 128'b01101100010111011011011100111001000000110101100100100111011000010100001100110110110111101011011010100010011101011110100101010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2778[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2778, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111110110101100100011000000100010111111011101000010101001000000111101100111111111101100101011100000100010010000010010011000; 
out2779 = 128'b11011000011101001000001110000000011010111000000110100011001010101101111110010100101011100001011010011100110010110001001101001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2779[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2779, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100011111001010000001011011100010111010011001100000111101000111011010101101110010101000110110110000001001001000010110001011; 
out2780 = 128'b00101011111100011110101010010000110011010100111100101101001100101101110000010010100111001010000111111001101001011100111000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2780[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2780, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010011000110010101111011000001101110111011011001000110000010111001111100100000110011100110101110111001001011111011100101001; 
out2781 = 128'b01110010010000101110001111100100000011010001101101001100100111010001001110111100101111011110011001010111010001000001011010111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2781[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2781, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011100000110011100011111100100111110111100000000101100110110001111100111101010110110101010000000100000110010110110101110000100; 
out2782 = 128'b01111100100111001001100111000110011010011011011110010101000000001100010110100111111001010001111101101011111110110010010010100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2782[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2782, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011101000101110010000101110100111001111111010100001010101100000000100000101101100100010110110010010001110101001110010100110; 
out2783 = 128'b01011001001110010111011100101000001001000111100011100111000101100101010000111000100011001000001000111110110000011101011111101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2783[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2783, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001101100010100111000111101000010100000100110011011111111100111011110010100101011000111111110011110111011111101111010000010100; 
out2784 = 128'b11100010110011101111110100101011011110011010011100011001000000000100100001100111000110001100010001010000010001011000001100110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2784[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2784, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011010110001001001011010111101010111101100111100111010000100111010000101111011010000011111000111101000101110100001100101110; 
out2785 = 128'b01000010011110111011101101101100010100100000100010100011111000111001000001111110100110100100111000001010000010110000011011001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2785[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2785, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111001110000010111000010100011001101000101100010001110100011001100011000100011110001000001011011010001100011100010100101101; 
out2786 = 128'b10011100001011010010010100100111001010100000011100110011100111010010001110110110100100000000011000001111010110111010000011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2786[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2786, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101101100001110001101010100001110101100110101000111011011110001100001100001100110001100110011111001010110101000100000010011; 
out2787 = 128'b01010100000011110000101001010101100110000011001100110101000101100010001100101100000101111001110000101010110001010100110011110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2787[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2787, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110010110111011010111110010110100100111011011111110111000101000111011110110000001100100000010011001111101001000001100110001; 
out2788 = 128'b01011111110111010111111001100101111011000111101010111001001101100000011000111010000001001000001010001000001110100000110010100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2788[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2788, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101101110000010111111000111011000110001101110111111000011101001000101111110110010001110101011000110001100001001100110110101; 
out2789 = 128'b10011111101010111000000001010000100000100101101100110111101100111111011000000110011010011001111111000010111010001000001010110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2789[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2789, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100101000100011001011001010111111100100111101100101010110110011110111100011100110001011000001100000110001100010110100111100; 
out2790 = 128'b11101011100110001100110111011001001010001001101010001010100100101001111010110011101011010101101000101101000000110110010100111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2790[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2790, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001001011001011010101001111101100100011110101111110111011110010011100110101111100000101011001011111011000010100010001000110; 
out2791 = 128'b11100110001011010101111111110010110110011100001110010010011011000010011001010011010001100001100111101110001110000101110010100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2791[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2791, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100110110100010101010111110010001100010010001001101001010101000101000010000001011011111111011000001110100010010101001100000; 
out2792 = 128'b01101010111011110000001111110011100001001000001111001100000110100111010010110101011100110111011100110100010001101000111110111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2792[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2792, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110111000110100011010001110101011101001001010110001111011011001100011010111010111010101001100011001001001000001100111000010; 
out2793 = 128'b00100110001010101010101011100000001100000010101011000100111001101101000001100110101010111010110101100100000010011010110010100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2793[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2793, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100100001011111000000101000111000001111011010111011100000010011100110110100010110000110000011000100100111100010111011010100; 
out2794 = 128'b11001100111110000111000010000100001101110011000110111010001101101110011101010101101101110110001110001101100010001111111111001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2794[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2794, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111011010001000001110010111111011010000111010110010010110010000111100111010000011010010001001001000011010110000111110101100; 
out2795 = 128'b00110100010011000011111010101110100010101101011010010011000001010100000100100000011000111111101000111111111000011001111011010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2795[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2795, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011100100101010010010100000101111001101110100100000100001110111101010000110111000100110111100110100010101111010001111110100; 
out2796 = 128'b01000111110000000101011000001001011111001101111111001101011111001101001010000010000011000001100101111101100110100011011100101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2796[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2796, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000110110101000110100100001101111010011100101111010110101001101101011100001001111110110010010001010110111000000011001100101; 
out2797 = 128'b11110001011101010101111010100110011001000101001011110000101011110111101100001011000011110100101000101111100100001101000000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2797[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2797, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101000110011011110011110000111001011111100100010110011110101001000001010000111000000010110000101011110000011000010010010100; 
out2798 = 128'b10100110000111100000011001111110010100111001100101101010100110000010110011101011111101101010100010011001110011101100001100011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2798[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2798, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000110111010111101011001101101111011100000100000101010000010111000100000111001101001101011110100011100001001000100001001101; 
out2799 = 128'b10101110110000110010111101000111100011001100010111010110110000111010100111111000111001001110001111101010101010001110011010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2799[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2799, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100000111010011000101010100010101101111101111011111000110101001110101001110111010110011001111101010101101010100001010101111; 
out2800 = 128'b11101111001000011010100001001100101001000011111011010000011110011000100011000010101001110100011000010111100011111111110001010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2800[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2800, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100000110110101010000011100010111100011000000011000111001010000000111001100010001001011101101101000010111100010101011001011; 
out2801 = 128'b01101001000010101011000100000011001011011100100000100100010111010111111010010001010100010110100001011010101011010010001001000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2801[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2801, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010111010100000100010001111001011101011110000111011000110000111101110101011011010100101001101101000101001100001000010110101; 
out2802 = 128'b01100101100001001110010100110111010011111101100100101001011000101010011111001011100101011101001001001111011100010110011010010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2802[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2802, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111010010011011010110001101000110001001100010010101110101010000100000100101001001110111001011001100010100010100010011011011; 
out2803 = 128'b11010010011011010110010111011101011000010000111101001000011110100111000110100001001101111111101100001111110111111000001011010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2803[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2803, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011100010100111101011010110110011000011101111001111100000110101100011101001101000001101101100110010111001010110101001111110; 
out2804 = 128'b01010001010000001001011000001010000101010101101111101010110101111000011100111000000011011110110001110111110010100001001001000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2804[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2804, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001100001010111001101110110111110111110010100101110100010011110111011111101100001011011010100001000001100110010011001010101; 
out2805 = 128'b00110011101110000000101101100000001100101000111111001000100110001111001011110111111111000011110000100110101000110111100101000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2805[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2805, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110101101111000000111000000110100100010110001000010100101110001111001111111101110000000110100111110111110011001111010110010; 
out2806 = 128'b10110111011100110100101000011101010010001010101000101010001111100010111111010010010111010101100010010101100110101010000110100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2806[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2806, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010110001100100001010000000111000011111110111110101111000010101001010111001001100001100010110101011101001110110011000000010; 
out2807 = 128'b11100010110100000110010101001000110100101010100101010100111101011101110000011001100111101000110000010100111101101111011010010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2807[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2807, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101011101010000110110101100101111000001111010000001111000100111101110111110000001111111101001110000101010110001111101001001; 
out2808 = 128'b11101000111000111010001000011010101100011001110010011110101001001000000111001001100111111010000001101001000111110111111011011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2808[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2808, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101011000111110110100010111101110000010100000111111011010110011100000111000110010010101010000011110010000011110001010110011; 
out2809 = 128'b10001100101100100011110111000000000100100001101011010111011100101100111011101111001001000001010001011010100110101011000110010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2809[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2809, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110110001111010011000110001101100011110000001011110001110110011010111011100000100001010000001010111000101010111111110100101; 
out2810 = 128'b01001011100010111100000111001110001100000000110011010010011010110111010001101010101101000101100111000111101110010000100000100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2810[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2810, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001110010110000111000000101101001111100111000001101001001000010110011001100110101100111100110111111001101100101111101101000; 
out2811 = 128'b10100010010101000101011100101111111100000110010010010111001001110100001011000000000100100001011011010100101000000010001000100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2811[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2811, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000111011111011100101001111001000101011111101100101101010110111111110100111001111100111101101101100011110011001001110011110; 
out2812 = 128'b00010000000010000010010110000110110011011010010111001010010110101010011100000111110001011100110100010000000111101000011100101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2812[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2812, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001100100000100010010010110010001000010110111001000001101000111010100011111111000010010110110011001011100101100100100111101; 
out2813 = 128'b01100101001011101001000100111001110010010011010101110101011011010010000000010000011000011001001111111011110001111101100010111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2813[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2813, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011000011011110011000000011101011010101011011101100011001001111100001110101001011000000101000110100100001000111001010010100; 
out2814 = 128'b10110101010101110110010101001110111111100100001111110010100000100110011101111001000101101110110110100000110010111101100100000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2814[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2814, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010011011001000101101011111101001010011010011110111110110111000000011000111001011111111011010001011100011010000100010110111; 
out2815 = 128'b00011001001011100101100010010011110000001110111111001010101110011001111101100001110010011110000110110000100001111010010010110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2815[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2815, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011001010101001010011110100100000011101001000011010111001000111001111110110110100100110000000010100011101000111110010111000; 
out2816 = 128'b00101001101110111110101001000110000101100100100101111011001100100110111111100101001001110111101001101011110100010000110110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2816[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2816, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111100110110101111101001101110101110000100011100100011111010110111101001011011110111000000101101000010101011011011010101010; 
out2817 = 128'b10101110101101100011100000110100001100011001011110001000011100100100011000111010011001001000011010000011101101010011101101111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2817[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2817, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101101100110011000010110011000001110101000000110001010111100001010111100100000101111000000001110110000111100000001000101110; 
out2818 = 128'b10101100101011100010010001011111011101000110000000011101000000000101111000010011111001111101001111011100100110101100010110111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2818[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2818, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111101111001010000100011101010100000100111011001000010110010010111100111100111010101001100101110010010110111011110010101010; 
out2819 = 128'b11001101000110111011001100000111100110101111000000111011111101101001100010011100111010000100001100000100111101000001100111101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2819[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2819, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001001010111010101000001000111110111111000001111111001010111111110110101111100111010011010000000001110100110000111100000011; 
out2820 = 128'b01000110101101100000011110101101110001100110010100111100111110001011101101110111111011001000001010101111111100100000001101001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2820[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2820, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101101000100001110001011011100001101111010001110100011100001000101001000100101011010110000100011000110001110001101010001100; 
out2821 = 128'b11010110101100000100000000011011011110000000101101000111001101011101000110111111110101111111010011100100000111000000000010010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2821[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2821, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100010101011010100001010011000110110011010011001001101111010011110110011100101110110100110011111100010100111001110010010110; 
out2822 = 128'b10110011101001010001000000000101001000100101000111000011100000111110101111001101111100111111000010001001000111011011101011111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2822[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2822, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010111010111110101111000000110101011100001010110100010011100111011010000111010110000010111001011000101011010000101111001010; 
out2823 = 128'b11110110001001101000110001010010000010010011010011100100101100100100111110010011111100101001101000001001010111001100001111111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2823[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2823, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110010101100010010100000010101011000110111110001011110101111010011001001000111000110010001000001001001000001100011111111011; 
out2824 = 128'b11011010110000110000000011100100010000010011110101101111110101110111001000111001110101100101110101010001101001101111101110110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2824[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2824, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001111010001010110000000111000010011110000011010000011100110000111101000011000111110101010010101100101001001111001111110011; 
out2825 = 128'b11101001001101001001001000001010011101010111000111001100011001100110011000011110000011011111011111000101001100110101111100000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2825[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2825, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101011011010110110001001000011110101000101111101101101111101110001110100111110111000001011011000000101011110010000001011010; 
out2826 = 128'b00001110011000011101101100000001010010110010100100100111111010010011000100001011111110110011001001000111110010100111111110101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2826[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2826, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101110000010011001110100001100110011001111100010011011101100110101011001001111101110100111110010010100111001110011010011011; 
out2827 = 128'b00001000110001011010101111010000100011000101000011100100001010000000011101011000000101001010010111100110110000100100011000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2827[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2827, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011101010101001110111000000110110110011110100010111101011001111110101000010101010100100101000000011000110111001110011100110; 
out2828 = 128'b10001110101110100100111101100010100011001101111011100101001000010101110001110111011110101101000000101010000111000000000101001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2828[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2828, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001010010110110001111111101110111110101010000010011101000001000010000001110010010110000111100011010010000100010001011000100; 
out2829 = 128'b10101000011000001111010000100011110011101001010011010110100011110111100110010100000010001100101100110110110110111001111011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2829[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2829, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010000101000011001111001110110111011001001110000010111101011011010011100100100001000111011000111010011100001111110101100000; 
out2830 = 128'b10111011000000011111010100101101111010000110111011010011011100100100010000111010001010100101110010101011010000000101010011001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2830[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2830, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111000110000110100010110110110101110110110000100000101001010011110101010010100000001110001101011110011100101010101010000101; 
out2831 = 128'b00110111001000000011001001100000111101111011011001001000010001110010011011011111111010001110110000010101101100111011110000101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2831[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2831, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101111111001010110010011010010011011000111000111001000100000010011000011110010111011111101100010101011011110000011100010101; 
out2832 = 128'b11011111100000001001011001001101111100100110000111100001001001100010110011111011001001111001111111000010111001110101101100111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2832[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2832, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000111001001111110111111101100001011110000011111111110111111110111110001111001111001100011100111001010011100110111010000000101; 
out2833 = 128'b11100101111101110010101011010110100010111011101000000010000011000111001100001011101000001111010000001010110001001000100001100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2833[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2833, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001000110101000110110000011110110100001110110001011011101010000011011101110101110100101101110001110111111001001100001101010; 
out2834 = 128'b01010101101011100111111010111011110010100010100001110011100100000001011000101000000000011010101011100010110110101010001000111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2834[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2834, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100000101111101000111000111101000010000111110001100000001001110011011010001001000000110110111110101001110101011011011110101; 
out2835 = 128'b00101011101100011010111111110111000101111010111111100110110010000110011100001010010001101001111100000001001000001011000011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2835[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2835, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100011100001111100111000010011001101110000000000000111010001010001111011100100100111010010011011111010100000000101011101100; 
out2836 = 128'b01000110110111101000101100001000111011101001110011100111111100010010101011010001110010011101111111100010110100001110011110100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2836[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2836, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100010110010100101001000110101001011100111100010100111001110001000101101111001101110100001001110101001001001000001010000011000; 
out2837 = 128'b01000011100000001110101011010001001011100101010011100001011010111000111011101111101100111111010111010100101000010100101011110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2837[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2837, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101011100110101001011000110110110011000110010000011110001101111100011110111010010101011100010000010010101110001001000110101; 
out2838 = 128'b00101011011010001001101000000011000111001100000000101001000100001110001001001001000110100010000001100010011001110100100101000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2838[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2838, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101001000010001111111001111011001000110011010101010101011110110000010100001111011110011100110011111100010010010111101111110; 
out2839 = 128'b11010110100110101011100000010100101001100100011001101100101100110101010011100010101011101111000101001001111010011110011011110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2839[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2839, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011110000111000011000100110100110110111011111110100110111110111010111001000001000000001011100011101111010010101110010111101; 
out2840 = 128'b11110111001000100101101101101010101001010110110010010101011100010011111101001011001011010110000000011000101101100101000011000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2840[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2840, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110000010010110001110000010110110110101101101000100000101011100001110101011011111110010001010011001010000001000111001000010; 
out2841 = 128'b01101100100011011101111100101000110100110110011101000111101110101111111001101001110110001001000100101111000101100011000110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2841[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2841, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011001111101001010111100110111010101001000111100001111110111100001100110001010101011001011001001110001000110100001011000110010; 
out2842 = 128'b00011001010110011111110000111011010111101100001110101001011111111001010110111111011100100111110000101110011111000010100001101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2842[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2842, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111011001101100001111111000000010001001010100011100010111000010011010011000011011100000101111010101111110100100001000101001; 
out2843 = 128'b10000011000011010101100010101010101110001100010010001000010010100001001101001111000101010100100100100001100000100110001111111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2843[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2843, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100100001010011010001011000011010110000101110000110011010011111110101101011001110110110110111010010111000110000010101111101; 
out2844 = 128'b10110101010111100101010100110111101111101001111111111000111001011100101110010000001111011011000111001011111011000011011111001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2844[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2844, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000110110011110110011111010110111011100011111100010011101100011010001001110101100100110101101111101000110111110011110101011; 
out2845 = 128'b10111010011101010010110111110010110010010110011010110010010000011010010011010011011001000010100001001000000101001101101111011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2845[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2845, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001110101010010010110000111011100010000011011010100101100101000001001010000101101110010101110110111000111010100111101010101; 
out2846 = 128'b10010111001101010110000100000111100010101011111010010001101010110000001010010101011111010000111101010110001110010100101110011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2846[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2846, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101101011001110100110101010000100100110101001100110101011000010001011110010100001101011100110010101000100010000001011111111; 
out2847 = 128'b11000110111101011110111010111101110100010010000011000110000110100101111001101000011101110000011000001001101100001001011100000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2847[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2847, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001100001001110100111111110011111101011100000110101100010110110011001010011100011000010010000110111010110100111100101000010; 
out2848 = 128'b01011110000110010111101101100100011001010000001011000110011000110010100010101111101000101111010010011001011000010111111110001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2848[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2848, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101001100100001110100010111100011110011101011101101111000010110100101111110110001111111011010100110101110101000110001000110; 
out2849 = 128'b00011000010001010100000001111101101110011111100111011100001110101001011100001111011000010010001110011001001110110100100010111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2849[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2849, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010011011010010101111101111101011000010001010001000111111111110011011000010101111001100010111111100101011100001000010001101; 
out2850 = 128'b01010011000100001000000011101111111100000101111011110011001100010110100110001001000000101010011011100000101100110000000001110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2850[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2850, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000110010000010010011011111101111001111001001110100111110111110100000011010000010011001111100101011000010110111011110000001; 
out2851 = 128'b00100111111001101110011101100100011111111000111000001110100101101100011000110111100100101100101001011011000001001111111011011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2851[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2851, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001100000001111110110101011110100010111100100110010111110000000111011111010000100010011010111101010111111111111000100010000; 
out2852 = 128'b11000111110111001101110101011011101011001101110010001011011111001100001000111000111001111111100100001110101010111101101001010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2852[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2852, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001111000101000000111011110101100110100100010010001011100101000001111001000011001110110000110110100101101101110111101110001; 
out2853 = 128'b11101001011010100001010110000110011000011111000000000100011110101111011000100011010000010011000010000110010001011010111011110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2853[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2853, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011101101111011111000011101010001101101100100101110011100011001101000000111000001000001011010111110100000010000000110001000; 
out2854 = 128'b00000101100000000111001001110110111110001110100100100101001110001110111100001111000000110001111010100000101000010111100100110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2854[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2854, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001101001010110101110001011011010100001011010100010000011000111001000011111110111010000110001100111101101010110011110000111; 
out2855 = 128'b10100100010110110110001000100000010100110101011000100100001100101011000110111011100110111101000010111010100100100100011011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2855[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2855, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001001100100000001111010001110000000001010101010001011111110101011100110011100100101011011001100010110100011111000000100110; 
out2856 = 128'b01001010101011100110100001110101001001010101001110011101111111110010011101110100110001110111001001010111001100000011111000100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2856[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2856, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001010101011011000000011011111001111100001011100101000110011100000101100001111010010010101010000110111001110001011111011111; 
out2857 = 128'b00010110011000110101111111111111010011111110100010010111111010001110000111011100011111000111101110001110100011000000010010010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2857[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2857, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111100101101000100101000100011110000100111100001001000101111001111000110011000100010101101110101100010110100001111010010101; 
out2858 = 128'b01110111011101111101000110111000010111100010001010101110100000011010111110110011010110011110100111010100010010100000010011011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2858[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2858, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110001100011111100010001011110111010010001001101100010100101101100001110111101100000000001010000011101101110110110000001110; 
out2859 = 128'b11111101000101100101000001011110101001011111011011011101001000101010101111111011010101001110011100001010010011001110100000110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2859[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2859, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011110101111101101001111111100111101110011101111101010101101100000001000110010100000000101000110010101101001011111101110100; 
out2860 = 128'b01000110000110100010101110011010010101000000110110000101101101100000110010111001110110011010001010010100110110001001101010010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2860[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2860, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010101110111010100100001010101111111001010100101110011001010110110010011110110101011110111100011001000100010000110011011001; 
out2861 = 128'b11111000110000000110110111101000011101110111110011111111100101011111001000111110110110111101111000001010111011110001111010010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2861[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2861, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111101100000111101000010011110001100001001000110111001000101110001111110001011111111001101001001001001000111001010101100111010; 
out2862 = 128'b01100110110001001000011101001101111100000001000101111011010011101000001000110011111110100010000001110101001110110111011100101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2862[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2862, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100001101001010110011000011101111110100111001010011101100000010101011101101000110100001000101101110100111101100011010111000; 
out2863 = 128'b01110011011011000100110011111111001000000000010110101000001000110100101101110000000011100100011000101011001110011110100011001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2863[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2863, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000111011111000110010110100001110011110011110010011110001110111100101101010010101011001010111111111011100110101010010000110000; 
out2864 = 128'b11101000100100000110111110000101111111111101101011101111110110110111010010100101001100000100101100101001010100001010000111111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2864[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2864, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111011101010111011110000010110101101100101100100000011100011110101001011010111101001001011011001110011110110110001000011111; 
out2865 = 128'b10011110101011000001111010100001010001001111010100111101011010101011010001111100111001100011010001010000001000010101101001111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2865[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2865, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100010001011111111000110111100000110010011100111010110000010000011101010100000101101011001111000010011010011101000011100111; 
out2866 = 128'b11101010011100100000010000011101101011111011011100010001001011010111000111000011011011001101011111110001110010101001010111101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2866[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2866, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000111110101010010010011001100010011000010111111001001000010101000100001000101011011000100001000100100111110011101011010111110; 
out2867 = 128'b10110101110010000111100001010000000000000011011000010011110110101010001110111011001100101011101111110000000010100110011011000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2867[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2867, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001001111000110100111110101100010111110001111101111011001010001110010000010000100001000011100100110111110011110011011000011; 
out2868 = 128'b10000100001101110010000111110000011010110101000111100111000011100100010101111101110011110101111111001000010010100000111010100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2868[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2868, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001010110110001111110110110010001111101111011101000101101001010001111000110101010010001000111110001010100011111011110100000; 
out2869 = 128'b10100101100101100101010100101010001100010010000111001110010110100110111101010111010000100111100110101101101011011010110110001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2869[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2869, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101011110100101011110011011001001010100010111001010001111000011011111000001011110001011111100110110010100001010010001110101; 
out2870 = 128'b11110010101111110100011110000011001100111101010001001000000110001100000111101001011110110111110111100001010011100010101100110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2870[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2870, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001000100001110100000001110010110001000000011100010011011000010010110010010000001001011111000101101100110010000001111111001; 
out2871 = 128'b10111010000111100011011000111111001110111111000010101010001010110100101101100100010111001101011101110110011101011111110001011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2871[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2871, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100101110111110100101111111001011110101111110101011001011110001000011100101110000001010000100110100011001011010000101011010; 
out2872 = 128'b10000010100001010000001001001000001111110011100001101100110111101111010101111101110100100101011001111100011111001011100101100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2872[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2872, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111001001101110001000100000011000000011111010000011101000101111000101101110111101001000010000110010100000000001011110100011; 
out2873 = 128'b00101101000110000011101010110010011111001000010111011000011011011000010110110010111110101011111011110001110000100011010011001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2873[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2873, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100100111010011110101000111111001010011100001001000011111110111110011110001110101001010000110110011000010011100010111110100; 
out2874 = 128'b01110111010100000001101111000000000011110001111011111001001010011000011001100110011011101011010110101000101101000101010101010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2874[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2874, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000110010110011010100110001010101001000001110101001000111010001001110111101110110011110111101000001010101011110001001001101; 
out2875 = 128'b10101001111100000010101011011101101011100100110010100011001000011000101001101010000101110011000101011001011011111100110001101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2875[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2875, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010000000111011011010011011111000011111001001100110110001111000111100100001101000001100010101111111101100101110000010110100; 
out2876 = 128'b10001101100111111110001110100010001100011100011111110110110100000001010100110100000011011110001100010011000111001010010011001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2876[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2876, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101111010010110011010101110101001100000001101011101000100111100011010111000111000111011110011101110011100111010010000011111; 
out2877 = 128'b10010111101101100010101010011100010010110001100010001011100110001100010000101111100100111111011110110110100001010101011111011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2877[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2877, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010111110010010110110111111110100000010111100000001010101101111111011001011010001101001100011001111110100010001111111001001; 
out2878 = 128'b01011101001000110101101010011100111100011001100100000011101100100001010111010011100100110010001010011111000110111101001101101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2878[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2878, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011100110001111100101110101001000100011100010011101010100011001110101100110011010111011011101011010010111000111111100100101; 
out2879 = 128'b10100101110011111000000101111001001001011011001001010001110000111001000101010000000111101101111101011110110000111010110101000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2879[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2879, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101000010000010111001101000011111010101011110111110000111010010000100100001000010000111011011000011000010110110111011110111; 
out2880 = 128'b11000101001000110100001100110110111011101101010101101100000100100011101111111111000001011001101100000101010000111111100011010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2880[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2880, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100110100001011100011100010111101110111111000010001100110000001101101110110101110101100101010001110101010000010100001101111; 
out2881 = 128'b10100011010111010100110010110011101101011011100010001101111010101110000000001111100010010001001010010101000011010001011001110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2881[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2881, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100001011101001101010111000100100100000100100011010111111010000010100001100111001001011001011011110110110101100001110110010111; 
out2882 = 128'b01001010111001010001001011111101000000000001100101010000010001111101010110111110111011101001100110101111110010010001011100101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2882[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2882, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110100001001100101101000111100101101001100011100101001100111011010011101111110111001101001001011100100101001010100010001101; 
out2883 = 128'b01001111110101010110010000011110000111111010010100010000100001000000101011001011000011111001100010000101101111111001101000011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2883[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2883, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010101100111100010101111010111000011001101010100000101000000011101110101011110101110110111000011001100000101001100011010000; 
out2884 = 128'b10111111101000110001000101000000101001010111110110101001110101110101101011100111001101001000110110101110001010011010000001111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2884[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2884, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000010101010001101010110110010111101010010110101010011010110001100101000000011101111011000001110100111001001010111100010101; 
out2885 = 128'b01100010101100110010111001101110011110100011101110101101100000110011111111110100101111011000110100000000111100101100001111011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2885[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2885, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010100000100010000100000011001100001100000101011111001001000000001000010110110010000110010010000001101101101111010101110010; 
out2886 = 128'b10011101110011111110110000011111101001101100001101111111000110001011001001110011101100001110110100000110101100111001100010011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2886[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2886, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001101000110011010001010001000011110101100010110010011011101000000000110010011111100000101110101000001000010110000011000001; 
out2887 = 128'b01000110001110101011001001111100011111101101111100000010000110100110001010001010110010110010010001101000111001001100111001001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2887[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2887, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111011111110110101000010000000000010101111100000110111111111101011100000100100101110110001010000111101011110011110110011100; 
out2888 = 128'b01100111110101001010110001001111100100001010011000101110000101111000111110110010010100110101010101001011100111001010000010110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2888[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2888, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011111111111010000100011110110101011001110100110100110111011001000111111010001001101001001000110001101001010001010011001001; 
out2889 = 128'b00011100100100011100111000011110101001101011110111110101001100100001101011011111101101000101000111110011011001110111010001110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2889[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2889, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001011000101111111010110110000001000010101101100000001111010011010011010100101011001000010111011011100010100100101111011100011; 
out2890 = 128'b00001000011000011000100110100101110001100100011110101011010000110001001111111101001001010010111110101000010111000010011010000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2890[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2890, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011110100010111001111010100111010011110101001100011101101010100000111000110011000101010110001110000011101100100000110010100; 
out2891 = 128'b01000010110011000010101100010110101111110011000010100100001111111111010100101110110011010011000001011011100011100110001011000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2891[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2891, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111011010101001000110010110101101000110010101011011010111001101010100111001110111111010010011101110001000101101011111000111; 
out2892 = 128'b00100110100000010100110001010001101010101111110101100100100010000001000001110101110111100000000010111000010110011101100110100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2892[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2892, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010100011100110110110100000010010000100100110101001010100101001000011110000001100110100111010100101111110101011001101010001; 
out2893 = 128'b01100110100100011010011110111010101001000010101100001100001001100101010100010011000111111011101101010010010010000000110001011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2893[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2893, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101110100000110111001110010011101110110110110000101001001011001110101010111000011000001100110000010101101011010011110110000; 
out2894 = 128'b10010100000101101100001001110001110100110001000110101101101100011001100010101000010101110001111000110011111101110100011110011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2894[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2894, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010010100000001001000000001111010010001011000100000011000101110010111011010000011001011011001110100000001000000101101101010; 
out2895 = 128'b11011010011111010100011110011010010111110011100000000101010100000010100101011101111000010101010110101010101001110010000100010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2895[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2895, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010101110111011100001010101110001001000000100101111001101001000100110100001011010010011111001001011011001110100001010110000; 
out2896 = 128'b11100110110100011001100111001001100001010101000101101011010010001010011011111110100010110101001100001110011101100111111011000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2896[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2896, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100100001111110101110101100110101000110010111000110000110101110001001001010111111001011100001101101010111000100011111011010; 
out2897 = 128'b00101011000000101100011110011110010010100001001000000001100110110010110011110111010110010000100010000000011001110010000100011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2897[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2897, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011111011011110100100010000110100001011011111100000001100010110100101100110100001111011111101011000001100111111001100110101; 
out2898 = 128'b01001101000101111101101011110101001001110011111100001110001110111111001100110001100000000100000111100100111101000110011110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2898[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2898, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010010000110011011111100111010111100001100111111010011111001011001010110100000010001010111000111110111000011001001101100011; 
out2899 = 128'b01100101100101111011111100110000100101100111101001011100001000101111011001110010010101001011001100101001100011100000010110110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2899[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2899, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001001101000001101101100000010000110001100000010000000011100110111101110111111001101100001101011111010101011100000110001000101; 
out2900 = 128'b10110001011100010100100111110011000001110001001001010001110001111000010101001000110101010111010000110000011101101110110000001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2900[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2900, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101001100011011011001011000100000000101011011000000010011101001011011010000100001001000000000111110111101001110111110011110; 
out2901 = 128'b11011110101001100101000100010011110000001000010100011011111100011110100101100011110011110011010111011101110010010110101110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2901[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2901, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111110010110000000001111100111110011100111011100110000101011111100111100000011011110101000100011001101111110000111110100110; 
out2902 = 128'b01100001111111100100001101011000010011000111111101001110000101101111001101110011011001110001101110001100000111000100110000011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2902[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2902, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101011001010011101101110010011010100010011110011011000100010101011100001111111101010010010010110001011010011001001001101010111; 
out2903 = 128'b00100010110111101111100110111000100010100011101110100000001111110110100110000001111100111111010000010010101011000111100101101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2903[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2903, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001010011011000110001011001000000010110100110001101111001010100000001100101010110110111110100000110011010001010110100111101011; 
out2904 = 128'b10111111011000100000111011000111001011010010110000110010000010001001111101100100010010110101110000010110011100010010110110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2904[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2904, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001100000101100000000000000110001010111101001101010101001000011101001110100010011001100000111000100001101101001100100100110; 
out2905 = 128'b11101100110111001001110000000011110111111000001010101110101111110010111100010011000010001101110111011111000001011000110110011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2905[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2905, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111111000000111110010101011100100000010010110000100000101001000011100111101101111111001100000101001001111110111101000000101; 
out2906 = 128'b10000100011110100110110001101001111100010000110100111000111101101011110100011000011101010100100011000100110111001111100111111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2906[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2906, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000100010001100011001001111100101011110100111011000110011001000001110110100100100010000100011100111111101100001101011001100; 
out2907 = 128'b00010110100100010111110011111001101111111110111010110010111110110000010100110010110011000111100011101001100101000110010000000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2907[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2907, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011101111001001101111000010110111000101110001100001011001101001101001101011111101000000000111100011100100001010010011001100; 
out2908 = 128'b00010011100111010010011011111110000111110011010000001011000111001110100000001001110101100111100110010101001001101011001001111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2908[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2908, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101000001100110100101000111011000001001111011011011100000010010111011111101010100010010101101001011010001011000111100010111; 
out2909 = 128'b11010010100010111100100001011010001111100000110011000010011101001100011110110001000111110000011001111001110001011011111000000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2909[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2909, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100010010000000100011111101000100000101000101101101001110111100100001000010111001011110000110001111100011011101101011000100; 
out2910 = 128'b11100111110000011110111101111000000111111101011010011101111110100011101101011001100000110110000010001010010010000001010101110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2910[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2910, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111111111001001011101011011001101100101011110000011111011111000001001111001100100000101000010110100011100010001011010100110; 
out2911 = 128'b01110110100101010111011110100010100110101000100100110101111011110110001001111111001111011101001011101111001001110101110001101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2911[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2911, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000011111011101011001001100010000110001101111010011000001110011010111011111110011010101000100110011010101010000101111010100; 
out2912 = 128'b01111111011101100010000101011001010100111101101001100101111100001000011101000110101110011001010111011011110010110000101111111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2912[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2912, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110101110010011011110010101000001011110110010101101000011010010000111010100001001001010101000001010010001011000011001000010; 
out2913 = 128'b01110000101001001111110011101011101000101000111100111111001010011110100100000101100101010101001000110010101010000011001000011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2913[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2913, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011011110011011101001010001110000100011101001001000110011101101100110011101101100111001111001110101001110111111010010010100; 
out2914 = 128'b11011111011100101000101000011111010111011010000001111000110100110001111011110011111000011101111001011110010111011110100010111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2914[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2914, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101010001010000010000011010101001001100000111011100000000110111110100101011111100011011010111101011110100110001111000001110; 
out2915 = 128'b11111111000100111111100100101111111100110111011111000000101001111010011100000000011001010111111001111101101011110110101001010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2915[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2915, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100100110001100010110011011000011000101101110110010111110101100111100111111010010011110111100001011101101101001100011110101; 
out2916 = 128'b10010000001110010000111001111110111111101100001111000111011100101110010001110101001001100000100100010110101001011011001111111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2916[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2916, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100001101011011010010011001010001110101110011110011111010000011110111111111110110010001000010001111001001010110100000110001; 
out2917 = 128'b01011000011001110101110010111100101000110010001110011100000001010110011011011011001011001111111100000110111111101001011100011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2917[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2917, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101010000101101100001001110101101101101010110110111011100111011100100101100100110001100100010100100110111001110110001100010; 
out2918 = 128'b01011110010010110011100100110010110100010100100000010111010011010000100101101010110000011101010011110101110000000000110000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2918[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2918, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001100111100100000110010100010111111101101011010001111100111111110010000011100010010000001101010011010110010110101111110100; 
out2919 = 128'b00011000010010101110111001110110011011100001110000000000001101011111010011110101000000000011000000000111000110110110101101111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2919[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2919, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001110100001111011000001100100100010100010101001111000001101100010110010011100100011100011010001111011011001000000011000011; 
out2920 = 128'b01001001001110000010100101010110101001110010111011101111110110000110110000010001010011011010101111111101111000001111111111000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2920[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2920, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001100001110010000010101010110111011011110101110111110111101110000111000101011011010000000011011001111011110110101001011101; 
out2921 = 128'b00001011010100101111001000010010111111000000001010000000000010110100100110001111010011101111100011011100111101110001011110101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2921[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2921, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010100101011101101001001010011001110010000100010111111110010001001000000100010110000110001010100100011111111010101011000101; 
out2922 = 128'b00111010100000011010001110111010000111001011111101001011100100010010001010011101001010100010110101101010100011101100100100001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2922[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2922, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001101000110111001010100111011000100010011101010011001011100111000011100001011101001111011100111000100000010001100010001100; 
out2923 = 128'b10001011111011100111001111100001011011100001000010001000010110101011100010000010110111001100000111010101011011100000111000011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2923[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2923, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101111111010001111111101110101010011011011001110000010000111000100110011111001100011001111101101011001011000111010100000101; 
out2924 = 128'b11101001000000111011011111101000011010101111110001010010100010100110010001011100000101000001001111011110001000101010011101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2924[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2924, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010110110100000011100011011110110011010000001011111111111000101111111010101010011100100011100010001110101010000000101000001; 
out2925 = 128'b00011000010111111110000010010110001111110110010101110100010011011100011010100110110000001001011001111100100010001010001100001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2925[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2925, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011010011101100111011001101100001111110001101111000111101011001111101000110001101110010100101010101111010111111010001001111; 
out2926 = 128'b11111001011011111100100111110100011010000111001111101100010010110011001000101011101111010010110010011010100110001110110101010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2926[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2926, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010001011111011000011000010100100000100010000110100001100001000000010111101010110000001000110011100110100111011011100100111; 
out2927 = 128'b00101000010110101100010001100100010110000110001010111110110100011101101010011001010101011000001111101001101111010111101010101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2927[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2927, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000011101110100110010001001000111001111000010101000111001110111011111010000100110111110111100000110110101001110100000001010; 
out2928 = 128'b01101110101111011111001001100101110100010011010100110001110100110110010010011010110011101100111110100011110101101010011011100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2928[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2928, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001100001111101011111100010000101100100101001101100111001111010101001011011111000111000101000100011111100010110100001000110; 
out2929 = 128'b01001100110011011010011011010100101010100001101001010001111111001110101001100001101110000101000110111100111010101100000110001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2929[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2929, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101100000101100100110010101011001101000000010001001101000010001000001001010110100110010100011010001101101000101000011001111; 
out2930 = 128'b00000011011001010001010101000110011111111010101101010001101000011010011000010100110000100111111101001000101110111100100111000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2930[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2930, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011101101001010000000010000100111111111000001001010000110101011100111001110111001110000111001001111100110100100011011011111; 
out2931 = 128'b01010110010100111111000100010101100101100000111010001001010001110101100000111110011010111110100101001000111100011101001100011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2931[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2931, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100001101110111100000010000001110011010111000011000000010011101101101110110010010100110010001011101000000001010010111101111000; 
out2932 = 128'b00000011001101110101101110001111000001000011010101100011100111010110101000110011100000100010101110101000011010110001001111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2932[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2932, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110111001011100000111011110011001000010010001001100101101111000110010001011110000011010101011011100100010100000111001010101; 
out2933 = 128'b10010011111010001101000101101110100110011100000100101000000100011010111010110110001110000110001011010110101010111001010100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2933[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2933, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001001001011011011000100010100011110010011000010001001110110010111010010100111011010010011100101101001010111011100110100010010; 
out2934 = 128'b11001101110100011111010111010100011101000010011110000010001100110111001101011010010100111110111111101001011100110010100100010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2934[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2934, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111110111101101001111001011011011110111111111000000011000010101111001000001110000111001101100010011011100000110101000100111; 
out2935 = 128'b11000111000011000001110011001011010110111011001110111110110111101100010100000111111000000111010100001000111010100101100100001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2935[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2935, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011000011110101111000000010110000000101010000111001011100110111001111010100010111110000101110001010110011010010110011000001; 
out2936 = 128'b00101010000111001100011100011001110011110000101111101100110011110000111011000110000110000001000011111101110111110001111101111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2936[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2936, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001111011011000011011100100011110001101111110101000110001010010110001111001010100000100111010011100101000100001011001100101011; 
out2937 = 128'b10010110000100111000100011111000111111000110110100111010011011011011010110110100111011101100010100111101100010101001111111001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2937[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2937, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010100111011111000100100010011101100011010000110101100110110000001001100011011110001011001000100110101011101110110001110110; 
out2938 = 128'b10100100101110101011100110101110001010011111110110000100100001010000001111111010100101111000101111011011000110110100001011010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2938[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2938, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100000011100101010010100010100101110011011001110000101001100001110101011010000101010101100101100000011010011011011100110100; 
out2939 = 128'b00001111111011110110010100001110111111100110100001110010000100001001011110001111011011001101011111001100101011100010111011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2939[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2939, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101011001101100010100100111000000100100011110101110100111111100110001011000111101100111111001001110100110111101011001100101; 
out2940 = 128'b10000110101101011101000001101001010001010111000111000010001001010111110001001110111111001000010010001110011000011111110010011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2940[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2940, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011011110011111101010110100100101010001001000101110100000011101100010001100010101110000010010000000100101110001101001001001; 
out2941 = 128'b11001000011110011101110100010100010000101001100111010100011011100111001101100100011101100100101110010000100110111110010010110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2941[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2941, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101100001001011001111100001010100101000111001011001001011110101111001101010111011010011111001000000100000111010111100010100; 
out2942 = 128'b01100101000000010110100100111000100001010001011110000100001001011110011101010000111000110110110111110000110000110111100000001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2942[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2942, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010100001010110011011000101010011000000101001100010001000111101111000100010111001010010001111001111100000101001110111010011; 
out2943 = 128'b01100001110011001110100001000000111001100111110011010010001000110110101101111111011001010110100001101011110001011010100011100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2943[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2943, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111101001110011010100001100110100000111101111001010000010111011100110111111010110010110100110110110000110110100101100000001; 
out2944 = 128'b10011010100111011001011000110111001101101101111001001101101001000101001010100101111010001101110111101100001010110001100100101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2944[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2944, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100100100101111101011100101010110001100011000000100100001100111010111011011111010011101110100010010111101001001001010101101; 
out2945 = 128'b01000001010111011011110101010010100111011001101000111001111100010101100011100100101001001000010000010000101000000111010010100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2945[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2945, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000011100000111011100101100111110010001110111001010101000010111100101011000001101010101101100010011110000010011001011001101; 
out2946 = 128'b10000010001110001011110101100111000000011000110100111000010001100101001111111000010001110101111010011010111010001101100111100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2946[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2946, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101000111111101010101011001111001011000110110010001110011101101100011011110000111011101101100101010000010101001000011101010; 
out2947 = 128'b00000010010101000100100001101001001111001000011101011011110101101000110001100110001001101000100110010001011110101110000111011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2947[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2947, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111110010001100000101100011101011010110110010100010011100010110111110100000100110110101000001101000010010010011111000010110; 
out2948 = 128'b11111001110111111010000000110000001101010110110001101000110001001000001101001010000111011111010010100001110101101001111101100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2948[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2948, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111011111110101111101100100001110011110011010111010011010100000001001111110100100111111111111101001110001110001001111001100; 
out2949 = 128'b10110100100010110000001001101000111010100111010000001111110110110001100100100011001101000000011000101100001001000111001111001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2949[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2949, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001010001010110101010000100011101001000001100101001010100011100111010110000101100101101110101111101010010011110110000010101; 
out2950 = 128'b00110010110001111101110011100111011110011111000001101100000111111101001010010011111111100010111010100100011000101101001001111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2950[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2950, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110110111001010101001110001001101001011110111011101011101000111101011001001110111100001110110101111111101111000001010011101; 
out2951 = 128'b00100001101001110000100000010010000011101011001111010001111111001111011001000100000110000001100011010010000111110111010101100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2951[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2951, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010111101111000001011001001110110011110100101100010101010000001101101010001100101110110101110100011001010001110100101010110; 
out2952 = 128'b10100010011010100011100000001110001100110110100000111001110110011001011110100110001010000101101101111011011111101001111100001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2952[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2952, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100010110100101001101011001101100011000000100011010000001110101011010100111110001100011010100110011001100101100111100100011; 
out2953 = 128'b01100001110001101000010001101110001010010101111011011001100001000011010111100011100010001010101000101001010100011111001100101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2953[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2953, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110010000011011011001001101110101011111110010011000000001101000101010000100100010001100001111101111101100110000000000100101; 
out2954 = 128'b01101101101000000010010101000100011011001101011111101001100100111101011010000101100100000100110101110110100001101001010111011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2954[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2954, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110001101001100001010110111001111010101001010001101100000000100001111010100011101111100100111011011100000001110011101011010; 
out2955 = 128'b10011000100101101000010110010011111000000101110111000100000001011101111000000011010010010111101011010110010101110001111000111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2955[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2955, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101100111100100010100010111110011011001001101001010010101001101100011101100100011010000100010110001100001001100101000001110; 
out2956 = 128'b00000101010010100010011000101101011100011010000101111011000101101101000100000000110110011101011011100011101101111111000100000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2956[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2956, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010010111111100110011010100101110001100000000000010001111001101110001101011000101000101100010101011011101001011100000011011; 
out2957 = 128'b11101100100011110001111101000110100001000010001111010010110111000001101011111010100111000011110010101001110001000001011010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2957[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2957, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111001001110010000001000010111100010010100000001001000101101101111001000000110110010001111100001010101010011100111110000000; 
out2958 = 128'b11110011110010001010110111010110111000101010011100010011011000010111011010100000101000101010110100101001110011111010001100111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2958[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2958, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011111101100011110010101000111100011001010010000111010101001010110101010001001101110110100100100100001110100110111011110101; 
out2959 = 128'b01101110110010100101101001011111011011101111111101100011111110010010001011000101010001011001011101010110011101001011100110100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2959[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2959, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011101001100000101100101111110100100001010000101100101111101011001101010010010110101101010110110111001110100001010101001000; 
out2960 = 128'b10011011100000010010110110110010010001110110011111010101000000110000000011110110000101000100111101100101100100011100111011010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2960[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2960, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001010100001100001011000110100100000000110111101101101111010100100111101001000100110000000110100110101000111100000000110000; 
out2961 = 128'b10001001101001101001001001111100001001010101000010111100011001111110000000100111010100000111001100100001101100001100011011010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2961[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2961, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011010110001100101110011011011001111100101011111111110101111100111110110010100110101010101000101100010110101001000001010010101; 
out2962 = 128'b10100111111000011010011111001001001010011110001000101101000001100111101101010100000001010011000111001011111011110110101101101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2962[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2962, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001100110100111001010100110000001111101010101010100000110100100100100000101111111101100100111001110011110101100100111110100; 
out2963 = 128'b11111011110101101101011000111110111000000011100001101101001110010000011000011000000111011101001101110011111000010010001000000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2963[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2963, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110100000000000011000010001001100111001000110110101110011100001101101011101000011111011101101111000100100011110000011010011; 
out2964 = 128'b10001000000000000010000111001011110011010110011111111001001010011001100000110101101000000101111111110000011100010110111101000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2964[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2964, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110100100111100001111100100111110111001001100110101000000011101110111100011010100010010000001011011001001011010000100011000; 
out2965 = 128'b10110001100100111111010001110110000101111111000010101100011001010101110111010100101101011000100111101000011101110010100110001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2965[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2965, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011001110001011010001110000111011010000111001010010000111101011101011010011110101000000110001000011011101111110011100011110; 
out2966 = 128'b10001100001111010011110011010101100101001100110010110011010010110011100010010110011011000001010100111001001100101101010000001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2966[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2966, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010011010000111100101100110111010001011100000111010101100110100110100110100001001101011111000110100111001001111011010010000100; 
out2967 = 128'b10101010110111000111001011011010001111100010101011111001100100000001111111101001011001000110101110011010101000000101001101001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2967[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2967, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001011011100010011000010111001000000101110111000000000110000111111111111110011000111011011110100010110111001001000101000111; 
out2968 = 128'b11010001110011110111010011000001011101110000010010110001011010111100001110100101000100100011011110101010011111111011001000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2968[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2968, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110010010010000101110101011101000110010101100111001001111011100000110101011011101100111010010100101000100110011110011001110; 
out2969 = 128'b00100001011101100111111000111101001001011010001011110101100010000111110101111110110011111110011110000101010001010010011101001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2969[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2969, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110110111000010110111010100100010001101100010110010011000000110000000001011001000011011011100000001010000111100010100110101; 
out2970 = 128'b10110111100011100101100110110110011101111101010101101111101011001101101110101111100110110110111111111011001101001101000000000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2970[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2970, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111111101110101010001100010001011000110010111001001111100101100000101000100111000001011010111110001001011110110000101100001; 
out2971 = 128'b11000111001110001100100000001110100101011011011101111111111101111011011110101110100111011110011011110101011011011100101110000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2971[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2971, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001100100010110011111101001101111110100100010110100011011011010001000001010011000011011011101001010011000000011101000000111; 
out2972 = 128'b01001110001001111000010111100110011000100001110011000011010000100011001110100010111010000001001111010100001101011010000110110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2972[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2972, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101100101011011110010001010001010010100111101000111110010011110011101111101000101001100101100000001111010000001111100011000; 
out2973 = 128'b00101011001011101101100010100100100011000001100101011111001000110001010001000100101100010011011000111100100101001110101101110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2973[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2973, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111111001110010110100010101111111010100100010111101101000001000000010101100111001011110011001110111100101011110000100101001; 
out2974 = 128'b01011101011100111100011011001001100110000111111111101100001000011101001001010110010000010001100101001100010011110100001101100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2974[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2974, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101000100010100100111110100011011011010010011100110100000111000011110100011101000000011000100001000010010010110010110100101; 
out2975 = 128'b00101000001001101111101000001011101001101101001001111100110110101001111001111100101111001101111101010111110010010011111111100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2975[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2975, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001110101010101001100000010001110011111111001111001101101100100010000001111100101011110011001101000001100101110000010010001; 
out2976 = 128'b10100101001011001011011011100101000000101001001010100110110010110101101001010011100100110111011001000101100010010101011000000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2976[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2976, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010000100101000100010110010000010000010101111011100010111010000001010100111011001101111010101011000111111000110110110000110; 
out2977 = 128'b01001011001000010010101000100100010011111110011100101100100000110100101010100100010010101001001110011010101001001001110101000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2977[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2977, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010001111110111100110011001000011111101111101111100000000110010100100101111100100101000100110001101000101011001001000101100011; 
out2978 = 128'b00101011110110101001111101010010010000101101100010100101001101100010001001100100110000000001010101110101000110001111110011000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2978[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2978, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111101010100011101100111011000000100111100101111110010000100111100011000110001101100010101111010010011010001100101010000001; 
out2979 = 128'b00100010001111111111001100011011101110110001111011001111100000110000011111010110011011100111001110111111001000100001110001011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2979[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2979, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001100000110001001010001010010001011100101101011010101000101110111100111111011101100111000111010011000011000000001010100110; 
out2980 = 128'b01010011111000100000111011000110110100100110110000000001011110001111001011011000011110011000111111011011101000110110010011101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2980[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2980, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111000010111011110101101001000010001111101001010110111100101011011010100110111000111100100010101100100110100110111001111100001; 
out2981 = 128'b01100001100101000111111001101100110110111000110011001011110100110111010011011110101111100110011011111100101001010111001000011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2981[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2981, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100010101001101011100000010001001100111000110111000100000001000110101000001101001111111100100111101000110011111011101111101; 
out2982 = 128'b10010000000101100001101001110011110000011000001011111010111011011001101111100110101100100100001100101100101111110101010011011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2982[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2982, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001111001101111000110111011110000100101101100001110011111100010101101001001011101100001011001011011111110000000100111101001; 
out2983 = 128'b01110000101111100000001101101110001001110100101010001110111110010000110110101001101010101100010001011110111011101000101001001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2983[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2983, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101010111100001100001111111010100111101000001011101110110000100000010011000010000001000101011100101001101101001100111110001; 
out2984 = 128'b11010000111101111000101000100000010001000100110001001000101101000001010100001110010110011010101110110100111011001010001110110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2984[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2984, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110110111001111111110100101101010111100100011111010010001110101101011010000111110000101011110110100000001101001110010001011; 
out2985 = 128'b01011000110000001011001011100010111110011110100111010110110000100110001000011000100100010110101000101111101000100101101011110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2985[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2985, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110011000001010010110110010101001111101110001000110011000001011011110101110111101111011110100110011110101010010000101111011; 
out2986 = 128'b11111010011100100101111110101011110100011000010100101111000110000111011100110001110101101001010000011010110001111100111001110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2986[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2986, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111000100001010000100111111101100110010111110100111001010011001111110110011101110011001010011110001110000011101001000111011; 
out2987 = 128'b10000000100010101010100100110010001001001011011011111010110010101000010110010101010000000111011111010001111111100010000000010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2987[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2987, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101111010011110110101001001100010101010110111100110100001111111000000001100011111110010110000110110001101111000011000011010; 
out2988 = 128'b10001100000111100100111011011101101110011111010001101001011111101100001011101011100110101010000000000100110110101100000001100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2988[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2988, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110000101010101001111000111001010000100111110101011011011001111100011010110110111101111001110001100111011010111011001011111; 
out2989 = 128'b00101100100101000000011010001100100101000101001001101000001111000100101110101011101011111000001000110010010100000101001110000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2989[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2989, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111111000001010101101111000110001000001101111111001000010101000000011111110101000110011100010000000100000110101000001100100; 
out2990 = 128'b00110010101000000001111110011100011110100011011110110110111010010101001101101110000110000101000011010111110111101011011111100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2990[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2990, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100100111100001011101101000001010000100111101010000001001000100000000111001110000010101010010101101001101100111010111100100; 
out2991 = 128'b10101000001110100000101111000101000010100000110001110011000000110011010000101000100011101100011000101001000010011101011010011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2991[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2991, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110011110100001000001000101101001101011010110110110010010010111101101101010101110011010001101100100011011010010011011011110; 
out2992 = 128'b10001101011110101100001101001100111000111010010011010110100010000000000011111111001010110100101001001110010011111100000000111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2992[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2992, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110100111011011110111100100101111000011000011011010110101101000001001101010001101111101000011111001100100010010000110010111; 
out2993 = 128'b11010010100010101111011010110101001000100001000010010001010111010110011110110011110110101010010100001000101111011111001101000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2993[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2993, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010010111001001001111000110011011001100110101000001000100001000011000111001100010001000011111010111011000101111111011010010; 
out2994 = 128'b01111000011111001011001011110100011001010110111110011010111101110101000111001000101000111010000000100001010000010100010010101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2994[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2994, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011100011010011001110100110000000010111010110010011010011110011000000000000011101111100110000111110010111001000100111011001111; 
out2995 = 128'b01001100100101100111010101001000101001001111100111101000111101100010000001110010011101011010000111111000000100100111000010110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2995[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2995, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111000011011000101000011110100000001010010000101110110001001110111010010001111011101010001111010110001110010100111110001101101; 
out2996 = 128'b00111111010010000011110010110011001110001111010100001101110111011001010111110001011111011101111110101001001110001110100010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2996[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2996, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010011100101111000010001000000010100110101110001000110001000100010001100101000101010101110101000101100010010101100111101110; 
out2997 = 128'b00001111000010111000010011111111011010110011001000101100000111110110011011110111000100111110001001010001011000110000001100110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2997[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2997, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110001010000001111100011001011001000010000111000101011010101000110100001101111011000000000011100100011111011110110100010001; 
out2998 = 128'b10101100001110100001111110111110110111111001001010000101101100101001101101000000010000001110011010001011101110011011000111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2998[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2998, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010011101000101100101011011100010101101101011011010101000010111000110001001111000110011010010100100101101001110000111011001; 
out2999 = 128'b00010001100101011101101110101000111010011101001010100010111110100100100100000011010011010100000000001101111100010100101101011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out2999[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out2999, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010111111100111011001001110001001111101011101101101011101111100100110110000100001010100111100100100111100100010001100111000; 
out3000 = 128'b01101000100100011111011101110110110101100111001001001101010001100001001110000001001010100111100011000001010001010111001110100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3000[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3000, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000110010010111100111111100011111010001001000111100101001001100000100001001110110010001101001100100101000000011100100000100; 
out3001 = 128'b00010111100010111011001000010110101011011010011010110011001110101111000011001101010000110111110100001011000110001001010101001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3001[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3001, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000000011101000111100010101100011000111001110100010101000100010000100111000100101010010111111011110001001010111101100111000; 
out3002 = 128'b01111000111001101000110010001010000010101101111100110101110011100100101110110101111110010010010000000011110010011101110010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3002[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3002, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100011000000101011110100010111100010011010010100100010010100000101000001111110001100110100001110111101100011010100011101100; 
out3003 = 128'b01100100110011111010011000100000111011000111110110010100011010111100110001001100011001010101010000101100001101100010001110111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3003[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3003, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110111101001111010000010110111010110001011000011110100001110010001111100001101010100000100100011100101100110000100010110000; 
out3004 = 128'b10001011111001011100000001110110011110001010001101010001000111011010011010100001111110010110101010001010000010001000011111100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3004[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3004, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001110111011110111110011011001001111001100011011111100010010100101100101010010101010000011001111110101110011001101001101101110; 
out3005 = 128'b11000000110011010100111100100110110000011110011111001000010110011000000110111101011000111000110110010000010101100010111110110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3005[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3005, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101100100010111101101100101001100011100110101001010000001011110000111010100110010111011101010100111110111110010110001101001; 
out3006 = 128'b00110111001111010111101000000000001001010111100111100110001100110001010001011001101110011110111010001100110100100000010000000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3006[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3006, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111000101000000101011101111111111011100001111011001101111111010001000110001011111111111011100010011110111110010101101010001; 
out3007 = 128'b00110010001100111101000100000111110100111111000001010110010000110110011111100101001111010011111100000011011010011001100110101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3007[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3007, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001001100110001001010110011001111100001100000000101111001000111111111100000100101111000111000001011101010101001101010011101; 
out3008 = 128'b10100111001110111111111101010100100111100010011111110100011010000111011101001001000011010110110101110011010011100001100111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3008[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3008, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100101110111100010001110100010010001110110010100111100001001100000001110000111010001011011110010011110000000100010111001000; 
out3009 = 128'b11110011111011110110011011011111101011001011010111000111001110000011010111010110111001111111010110110100101011010000111111011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3009[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3009, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111101111011001111001010011000011110011011111110011100111001100010000110111100011001101111010110100101111011100111010000101; 
out3010 = 128'b01011110001001011111101110011110111111100011110110000101000000011001100011010100001001000011010000001100000100001000011010100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3010[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3010, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010000011111011011101111100100001000010011110111011101100100110100001001101010101010100000010000001000000110110101001010110; 
out3011 = 128'b01101101100111111011001100011111001101010100001100101011011100001001101101010010110001111011110001000111001110110000011100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3011[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3011, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000111101111010110001011000110110011011110001010011110111011110000100001110101100010000001100111001011111010111000110001110; 
out3012 = 128'b00001100111011000100011110111111100000100001011001000100101000110000100011101011110100100011000100000111011101001111110111110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3012[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3012, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111110101100100000010110110001111100101100101101000010001000010011101010010111111101011100010000110001111100011000000000001; 
out3013 = 128'b10011000101011111110111111110000110011101001110000001011100011011100010110011110111110110011111111001111001001000111111001001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3013[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3013, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110100101110011111000110111011111011011001001110100000001101001111010110110100101101001111010101111110111000010101011101001; 
out3014 = 128'b10100001000011011010011110101101010110110100001000010000000100111010001100001001101100001000101010011110111011011011000001001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3014[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3014, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101011101011001000001000000000010010101011101111111011101110101011001001000000100100100000000110000100000111010011100001100; 
out3015 = 128'b01110010101110000101010110101001001101110011100110110011111101100101000101111000011110110010101110111100000010010011101101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3015[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3015, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111000110001101011011110111000110000001011000001100010000001001101111110100100111010110101011110101110111011000111101101001; 
out3016 = 128'b11101101100011110111011111001010111010110100011101111110100000100001110011011011000000100111100100011100101110110110101111110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3016[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3016, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100011010001100101101000100111010101010000011111101101101011100110111011101101011010000111110010100010011101000001001010001; 
out3017 = 128'b10101101000100011001101001100010001011001000110101101110000110110011000001111000001111001101000100110100100101010100101011011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3017[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3017, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001000001100100110101011010001000011111111010110101001001011110000100101011111111010110000101111111110110100110001001111100; 
out3018 = 128'b01001101010011010010000001101011001011110111111001110110011101100000100010000000111000111011100111010110011010101000000000100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3018[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3018, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010111111111001011001101110110001001101110101010101100111101001110111101110101000100110000111001001100100011000001010100100; 
out3019 = 128'b01100101100111001101111010100110110011010111101001100101011111010111011011001011000001100110000110000000111011111010101001101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3019[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3019, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100001110100011010100111110110010000001110110110100100001100100010111110001011011010110010111111100110111001101010100011001; 
out3020 = 128'b00100111010010010100101011111110101100001110011110111010100001100011000001011010010001000111010110010101001111010010101100101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3020[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3020, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111011110110010101110000110001001110001011001011011011010111100000110011011101001001011011111010101000101111110110101101010; 
out3021 = 128'b00001001000111100100101100000110000010010001011000101001101111000001101111101101011110111110110110110000001110111001111110000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3021[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3021, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111001011010011110011100000011101110001100010010000110100101111101011010010110110101010111110100011010010111010010101111011; 
out3022 = 128'b10110000110101110011110101001010111100000110011100110100101100000110101000010000101010011001100100110001010000100111101011010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3022[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3022, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100000110011111001001011101101001001010010010001000111011110100001001011100010010111101111000111001111100011000001010010001; 
out3023 = 128'b10001011010101011110111001001101001100010011100100011011110000011001001011101001000000100101100011101010000001100101111110110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3023[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3023, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111001001010100001100101111101110011011110110011001010110010111100101111110100001111000110001001100110000000101010010101000101; 
out3024 = 128'b11100011000000001010001101010010110010000001000110001101010000011110011110001110001010110010000001111010010011000011100111111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3024[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3024, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010010000101100010011110001000010100111001001001000000110000100011110111101011001110001110000100100111100101101001001100001; 
out3025 = 128'b11010000101000001000101101111001000100111001101111001110111111010001101000010010101110110011011000011010111001101000111000110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3025[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3025, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000111100011111111110001010011011101100101000110111011010101010100010001011010111100101111110001000110111110111110101001001001; 
out3026 = 128'b11111101000000111010111011000001000101011010001001000010010000010000100100000110010001010000000001101010100101110110000000010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3026[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3026, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101110010111010101101000010011101100111010010100110101011100101110101011101111000101000010111101011111010000101101010000001; 
out3027 = 128'b01000111001111000001111111110111100101110001001111111011101110001100101010011111001000110001110001110001100000001000110001100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3027[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3027, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100100011010000011100001000001011001100101100000000000000011001001011011100110101110111100111011101111011001111101100010110; 
out3028 = 128'b11110101101011110111011101001110010100001111011000000100111000111010101001010001011111001001101111110010111001110010100101000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3028[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3028, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110000010100111010100010011111100011101001111111111001011001110000110011110110000000100010101010010010100001110011110101111; 
out3029 = 128'b00111001000011001110101100101010111110111011010001001110110000001100000000000011011011101110100000011011010101000001111010100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3029[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3029, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111111001101000001001011110101011110010110010001111111000111010111010011110101000010001110110110010010111110110000111001000; 
out3030 = 128'b01001110011101010010100111111101011111000111000100001101010010100110010101100000110011001111100001000111100011001011010110110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3030[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3030, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000110001101110010011111111110110001110110110110010101010101110101010101111001000111100011100000110000110111000001110110010; 
out3031 = 128'b00100001111001000010100110101010110100111000100011001001011101111000000010010010111111000100111000000110001101011101001010001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3031[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3031, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111010110101100111001001011001111110100000111110011111101011010101111101110111011010111000110111001110110000001100000010101; 
out3032 = 128'b00011000000110001001101110101001000011101001111101101100111010101000110100111000010111100010111111101010101100100101000011100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3032[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3032, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001011110000110001011111011111010000101100110111001110110110010111100010001100001111101110111000110011101110011000110010101; 
out3033 = 128'b00010101011110110001010001001111011100110111011101001111010101111010110110111110001100011010101000110100000100101101100111011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3033[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3033, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100001111000011101101111110000001000011100001111111011000100011010001010111111011110101000111111110101100001001001111010110; 
out3034 = 128'b11111001010101101011011011010100000010111011101100001001101010011011000001110100110001110010001001111001000110000011011100110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3034[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3034, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001010111000100110100110010100111000101100111100000000000111100010100101100011000101100001101111110011101110110101100000000; 
out3035 = 128'b00100110011100100010101011101111000111010110000100110110011111010111111111101101111100011011001000101010011001110010010100110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3035[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3035, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111001001110000010101100011110101000001100000011101000010110101100000110001010001101010011000110010010010101110001010000111; 
out3036 = 128'b11010000011111100110100011111010011110010001111011011101100011000011010001101001111010001101000111100110101010001111000111111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3036[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3036, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100101111111010011101110011101001000100010110100111100111101101110110001010000110111011010001101100000001110011000011010111; 
out3037 = 128'b11101001001010011111001110100100011111010110100000001000110111001010101011010000000111001010110110000100011110101110001101100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3037[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3037, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111101110010001101011001111110110110101100010100000111100001000010001101011100000000011000111011010010111000011000010101100111; 
out3038 = 128'b11000111000101011111101101010000000100101100011100101101000101010110100000101101000010001000111100011101110110110101000000011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3038[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3038, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110100100110101001011110011110010000010001001110100000001110000110101101111100010100010100010001111101001100111110011110000; 
out3039 = 128'b00001110000110011001000101100011011110000111000010111010100001100101010010111110011110110110001111001101010100101101011011111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3039[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3039, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101110010001111101100000000111000010111100111111101111100101010111110100010110100001101000110001100111111111110110010110000; 
out3040 = 128'b11101110101011001111101001110001100000001001110011100010101100010011110110101000010110010100010111100110111000000011001110110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3040[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3040, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001001000110100001010001111000100101100101010011001101001111111000000110011000000001111011110010110001110010010010011000110; 
out3041 = 128'b11000101111010010110101110111110011000001011011111010001001110100011000110110000100110110101011110011010001110010000100010010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3041[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3041, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111001111110001101000000111100100100100101011001100111010111111100110010111000101001111010101000000010100111001011010011001; 
out3042 = 128'b00001000110010000101101000101011010110010001100000110100011100000101010011100011100001111000000110101001000010010010010011110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3042[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3042, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111010010010001110110111000000011011111001111001110011011001000001001000011000010010000110110010000100100010000100101100110; 
out3043 = 128'b00010111011110111101100001001001000010110010010100001001010011101111100100101101110010100010100011101000110001100101111101001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3043[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3043, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111000000010110010110001001110110000110000001101110001000101101100001101100010001000010010111100011100000010111001110110001; 
out3044 = 128'b10110001101000101111000001110101000101011010010011100001001111111101111010110011011111011000111001110010100010110110111100101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3044[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3044, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000111010100000100100111001101001000011000110100000001001011011001001000010011101011110011111100110111111001111100110001100; 
out3045 = 128'b00001110010001011111100110010111000010111100101111110010011110010110001001101001011101111000111111001100110101001110000101110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3045[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3045, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101110110001010110111100000011011110000101101101011010111011100010101010011111000001000000010110010101001110001001010011100; 
out3046 = 128'b01011011001101111110101100011010101011010011010011010000010011100100001011110101110010000010110101101000000110011110011101110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3046[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3046, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111110010000011010001100000000001101011100010001111011011010001111011011001011101011110100010110110111101011001010111001011; 
out3047 = 128'b10100100001101010011101101010100010011100101101010010110101000111001100001010000001110111010111001010101101100110110001001000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3047[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3047, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101101001101101000001010110110011101101101000100010101001111010010010001001000000000110010011101100100000110001101110001011; 
out3048 = 128'b01011110100110100011101100110010111000110000101100100110111100110100111100011011001101011000101000111010111000001101110101101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3048[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3048, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000100110110011001011000111000110010100111001111000010111001000100011000111100000111101110111011101101100001011100110101000; 
out3049 = 128'b01001011110100001001101100101110100101111000110001111111011011011101101100111011010100100000110001101001110111001111100110101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3049[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3049, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011001001101101111001000011100011010011110011011101011110011100111001011101110111100110101010011011111100001001111101010011; 
out3050 = 128'b10101111000100011000010111011000000111001110100110000010000101100001101000010100001000101000100011111100100110111000001111001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3050[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3050, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010011000111010110101100110000110110001011010010011101000100001110100110101101010001100010111110001010010010000000111111101011; 
out3051 = 128'b11001101000001101001100000000011000000111000111001001000001101111110000001000111111000100010010101001000110101000000111010110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3051[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3051, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000110010100101001010111110001101001000001100110000110100100010011100001001000110010101111001100011100110110101010110000110; 
out3052 = 128'b11101101110100111011000010011000101000011010101010111100110010001111000110010110011110111000010100100010010011000100001001000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3052[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3052, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001111101010110010011110010100001011011110110000101110010010111101100010100110111100000110010111100000110001101010110000011; 
out3053 = 128'b11101001001001111111000000001100000001000101100011001110110011100101101101000111101110011000010101101010110101000011110100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3053[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3053, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011101111000111010010001110011111001001100001010110110100101000000011010000110000100101111001110011111101000010101110011100; 
out3054 = 128'b11000110001010110110001010001110010000001000100110110111110101001010001110100110000100111101100011001000100000100011000100100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3054[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3054, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100101001011101000101111110010011000010010001101111101000010001010000110100011100110111101011110000001101010000010001000000; 
out3055 = 128'b10011110011101000011110101111101110001100001101111101111100001001001001111011111000111111110101100111101100000000010111111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3055[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3055, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101011100101011111111101000101111100011001001001011101000101100100000001100000010100110011000111100100101110000111100010000; 
out3056 = 128'b01111101111101001011111001011001110110110111111010101001010101011110011111000111000101010110110111011100000110100110101100101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3056[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3056, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110011111110110011010001111011111100000111011010011111101111011011110011111000100110011101111110001010000001101101111101101; 
out3057 = 128'b01001010100010110110110111000111001110000111111000000001110110010010111111100001100111101000001101010101100000000011110111100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3057[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3057, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111001010010111001100000111011000101000011100011011000000101000111110001111000110100110010011111010101111011001111100000000; 
out3058 = 128'b10100011100100001000001111001101010001000000011100010111110011111001000010111000010100110100010110101100111111001101111001010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3058[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3058, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101010001111001111111010100100001101011111010101100010100101110010111000111110100000100110001101100000101010110111100100000100; 
out3059 = 128'b10101110011101111100010010110111000110101001000101101000000011111110001110100111000011100101110001000011111100001110001000110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3059[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3059, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010000000111000101111000110000100101010010100110100010001011010011100001100000010110111100010011110100001101100100010100010; 
out3060 = 128'b01101110101111010101001001000110100010010010001110001011000101100110100010011111001000010111000111010001101111011111110010110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3060[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3060, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100001110101010111011001000000010100110010110011011101001111110100001000000000000100011101011110001011110100110011000011111; 
out3061 = 128'b11111000100100000101111110100010110000110011101011101100011010110110001011110101010011010110100111101000001101111110010101000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3061[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3061, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011111111101001011011010100011111111101011111011011001110011000110101111011010110010110011101000000001011011101101111000110011; 
out3062 = 128'b10000000110100100001011011101110011010010100001000011111011011011110110100110000110001100100101000011001010001101010100111100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3062[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3062, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010010101101011011001101100011100110000001000001000001100100101111010111000111101000100001111111110010110101001101111111110; 
out3063 = 128'b11000011110000100010111110001000010110100010010100000110011000001111101100101001010110001001111001110101100101100110100110010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3063[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3063, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001010101011110100100110110110000101110111011101101011001011101001001000010000110001100000000000110100011000001010011010100; 
out3064 = 128'b10100000000110110001011010010111111100001101001011110111110011100000110111101010010100010110010010000010011100000101000111011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3064[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3064, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100011010111110001001100010110111011010010000101110000110010101110010111110011101011111001001100110110000101110110100010011; 
out3065 = 128'b01110101111001111110100010010011010011001011101110001100100111010111101010101100101010100111100001011100111110111110000010000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3065[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3065, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101010100010001001101000111001100101010010010001001000101101001101110111001000010010001100010010111000111111111101000001101; 
out3066 = 128'b10011010111011001011001100010101010010001101000100011011111011011100101000011011100010101001101010101010010100111000010101111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3066[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3066, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100000010000011101111100110100011000110011110110001010000111111111101100111101101100111000001010011000001010101010011001111; 
out3067 = 128'b00001100001111100101000101111010010111010100110110110001101001111010001000000001000100010000110110100111100110010100101000010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3067[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3067, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101001011111011011010011011001111011101001001101101101001000100110110000101001001011001100000000110100000001111111011001100; 
out3068 = 128'b11110000100000000001101000000010111010010011100001111111101001010001111000111001010011110001110010000000110010010101101010011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3068[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3068, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001010111100111011001000111110010100010010001101110111010111111100010010000111010010100101101100010110001000100010011101000010; 
out3069 = 128'b01000101101110100110100011101011111101111000001100000001001001101011110111001110001101111100011101111010101111001011100101101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3069[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3069, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110101010110100110111010010001000011100110100011111011110111010001011000000001111000110101011111010111001110101011101010000; 
out3070 = 128'b00000100010110001110111011011110110100110101111110110001101011011010010110011010110100011011011110011000010001100111000110100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3070[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3070, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000110011000000001011101101001001100100010111001101000110100000011001011100010010100110101010111010100011010110010000101100; 
out3071 = 128'b11011100111101011001101101000001011101100110000100101000011100010100010010001001010100010011010010000101011000010110110011111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3071[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3071, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110100110100001011001110011000111110110101110100011101100010110000010111101101100111110001011100011000101110011110100111010; 
out3072 = 128'b10010010010011010000000010111010111101010010101000101111000100101010110000000010101000100010011011110000101111011111011101001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3072[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3072, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000010110100000111101000000110011000011100100000101000001011111111011110101110000011001110100011110000010100000000100110000; 
out3073 = 128'b10001011010100110100100110001110010111101110110011111101110101000110111111000101011110001011011111110100011101000000111111110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3073[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3073, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010000101010011001011011101001101011001101100101110011110101100010010101010101000001100111110011011001000001011010111011011; 
out3074 = 128'b01111000101110110100000110001110011010100100111101101011000110001001100111111110111010111111000001010000111001001001001000010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3074[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3074, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101110110000000111110011110010000101001101111110111001011110001011010000100110100111111000100100010110010111000001100111011; 
out3075 = 128'b10001011011001100011000111000100101101100001001101010100101000101010110001101011000000111001100010110100011010011101001110110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3075[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3075, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000010101111001011010010000101010100000100111100010100001100010110000110001001001011110001110111101100001100110011001101011; 
out3076 = 128'b11001001011101001110110110110101000001000110110111000000010011110100100111100101010000000001010100110110010000010101101100101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3076[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3076, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001001101011000001000011000010100000010110101100111101010010111110100000101100110101001110111111010010010000010011110000101; 
out3077 = 128'b11110100001010010111111010100110001100001000100111100101001110111000100010111100001001011010011010110111101100000010110101011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3077[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3077, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011111001001000010001100100011110011011101110000100011101011011000100001010111011101000010100000100000110111111000011001100011; 
out3078 = 128'b10111010111101101001101011000111010011100111100010101101110110001001101001000010101111010100011010101001001011000011010010001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3078[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3078, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010000010000000011100110001101111100100111100000010101110100001010100101100001010011000001111010011110101111000001001101110; 
out3079 = 128'b00101000011001101011010010000011100001111001000101010110010101101010010011100000110110000001011100000110011000110000100010001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3079[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3079, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100011011001010010100000001001111101011110111110110111101110100001110000110011010110111000000110111101001111101001000000100; 
out3080 = 128'b01011011101111000111101001000100100001100110111110001101111111011001100110000011110010011100000100111100011000100010111010110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3080[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3080, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001010010011011001101000100100111110010100011011011010110010011001010000010100001111011001000100000100010010010010010110010; 
out3081 = 128'b00110101000111111011001000110110001111101100000010000000000100101101111100100000111100000011010111100011010001110010101110110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3081[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3081, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011101010001110111100111100001100001011110101111011101001101111001011101111101100110001100100000101000010101010010000110001; 
out3082 = 128'b01010110011011111111001110000011101111100110001011000101100101000001001010101110000000110010011010110110111010110101011100110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3082[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3082, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001110101001001110100000010101001000011111100011011000001000000011110001101011110001110011100101010110110001100010110010010; 
out3083 = 128'b11010010000100111101101001100000001000001010010111010101101111000111001000000001111001101100110001110100101111000101000101000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3083[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3083, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000010110101000000011000001010111011001001101000100111000111100110010110101110000001110011000100101101000000010101011010101; 
out3084 = 128'b11111100101111011001001000010110001001101110110000001100111010010101111110100101011101011101011000000000100001101001001110010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3084[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3084, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110001001000000100011000111100101011011001100011110001001010100011100010010110001000100001001110010000011110111101010000110; 
out3085 = 128'b11100111010001001011000001110110000010110001011010010010001010011010000001011010000001110001101110100111011110001111011111100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3085[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3085, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001001111111101011100011111010010001110101111101111001011111110010010010000111010010101111000001110111101010010011110111000; 
out3086 = 128'b01011010010011000000101011000101001111100011110101001011000100000010110111001010010101000111111000001010100000110011111001101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3086[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3086, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101101000101101100100100101011110100010010110111111100011010010011101110111001001111110100110000000101101110101101110111111000; 
out3087 = 128'b01010100101110010100110000010111110110111101110111101000010000101100011101101110100010001010011111001111001100111101010010110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3087[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3087, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010010010110000110110101111111011101010011111001100110011111101000111001001111100000110000000001100010011010000111001011110; 
out3088 = 128'b01010111000010001011000100010000100000000111011001111101101011011000111011100110000101100110001000101011100001100110110101101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3088[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3088, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001010110111111110101000000011100100001010000001011001111101101111000000001001000011010101110111101011011100011011111011001100; 
out3089 = 128'b01000001100000110000010000011011011101001110011110100101001111000111110100001100001001000101000001100011011011011011001101000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3089[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3089, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001011001001110001101110001010000101010001011101000101011110110101001001101111101011101010110110101011000011011110100101010; 
out3090 = 128'b10111101101101001110101111110100000010000011110001000000111111111011000010100101100000010010010010000010011010100011011111111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3090[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3090, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011011100111011100100101010011101111110000001100111110010000011110100101000000101011110010010101010010111000001111011001000; 
out3091 = 128'b10101010111010010101111101010100101111000100111001110110001000010000110111100111111011100100011010100000000111111011111101010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3091[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3091, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100010000010011111001111000111000110000001110011010110100011110001101001100011111001011101100000000011101011000111010101010; 
out3092 = 128'b00011010011111000110110001101010001010100111001101110010000110010101110111001011011011100111011100010100100101111101101111001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3092[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3092, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000010011010110010000110010100001111111000100100001111010111000111100100110100110011101111000101111010100010110010010011110; 
out3093 = 128'b01101100011100101010000011001010110011100011100100100111011001010110100001110101110100000011100111111000111111001110001100110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3093[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3093, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000111110111000001000100001100111111100110011101011111111101101111110010100111011110111110001010010110101000011001100101001; 
out3094 = 128'b11110010100000110100110100010111101001100111010100100100000010100001001100110101010110101111101010011001010010101000110001100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3094[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3094, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000011001110101101000100110100101111010110110101111001001001000000000010010101011101101010010111101111101111100110001011100; 
out3095 = 128'b01000010001001000011000000100000010001100001110000011001101101011000101010110101010110000101101010011101100100100010000101111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3095[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3095, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100101011111110001010000100000010000000011000001110011111110100010001101111111100101111011110110100111001011110000011010011101; 
out3096 = 128'b01010101101101010101000011001100010000000100100010001110101111111011111010010101101110101101011000111100110101000110010010110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3096[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3096, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100110100010100100100001110010101011100110110110110001110000111100010001110000011000001000000011110001010010101100000100110; 
out3097 = 128'b10011110110011101001011010110000101101001110010100100111111010110010100100111100000011110011010100011110010010011111111100101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3097[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3097, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101011110100101000100000111111010101100011101100101000001100110011101111001000100001100111110001000111000110010001110100000110; 
out3098 = 128'b11101111010000011000101111110000010111111110110011101101001000110110110101110011100111001100111101001001100010110100011111100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3098[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3098, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100111010011001101111000011100010000110101010110010100000110000010110010101010000111101101010111010010000010011101110001111; 
out3099 = 128'b00110101011110011001011111100111010111110100101011100101010101010001001100000001000111110001111010010010101011100011001101101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3099[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3099, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011000001010001111101001001001001000100011101011110100111001001011010110101100111011000001000100000111100100101100100010000; 
out3100 = 128'b10111011010001110010011001100110011100101000010010001110000110111100100011011000011011001100000000000001101000100100001101001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3100[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3100, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110101000100001111101110101000001100011000011010101101101101100011111000011001011000110100100100010001001000000000001011001; 
out3101 = 128'b00110010001000010101110100110101000000100011111101010110110010100011000100001100010001011100011010111100110111110100010111000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3101[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3101, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001011000111111101101110011010001100101110110101011100011110001111000011110011011100010010111011101011010010001100010111001; 
out3102 = 128'b11111011001000000110000110010111001000011111101010001101010000001111100011100111001001111001111001010010010000101100001101110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3102[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3102, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000000010010001011100101000111000011011010000010111101111001011111000101100010101111011101011000010001010111111000011010000; 
out3103 = 128'b11011011000001100100100001111010110000100001111100101110010110011001001100011000100101111000010110011101101101000111111011100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3103[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3103, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011111100111111011110100110001000000101000100010111100011101100101011010001011101011101011001010110001101101001101101110001; 
out3104 = 128'b11101111011011000100110111101000101011110100001010000101110001000111101000000011011001010110001001101010110101001011010111100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3104[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3104, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111000100111001011101001000100101100010101100111100110110111101010000100111111011000100101011001111100100111001100101100110101; 
out3105 = 128'b11010010010101000000111111100111111101010011011110111010010110110000001001001111101110100010011100011111100000001101111111011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3105[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3105, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001001010110101111010010110000100011111101101110110010110011100111101101110110011101111110110001101111100001010011001111001; 
out3106 = 128'b01110101011101101110000000000110000101011111100011011011110111010011101101111100011010010100001111101111000010000000000001001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3106[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3106, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111101001100110101100010101110010000101000011110010010011111100100101001001100011111011011100101000111011111111100011101011; 
out3107 = 128'b11011111101101011110000111001111111111010100010110001011101000110011111111010110011001000100101000000100000010100001001010010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3107[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3107, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100000110110011100001000010010111010111010011110010111001101101100000000101000011100111110001100010011011000011101011111111; 
out3108 = 128'b01101011110111101110100010001001100111011111111110001101100101011011100110100111101011111000011111101111001011010110111111110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3108[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3108, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111010110010001101101111100100100101110000100011111001100100000110100010000100000101110001001000000010101111100101100000101; 
out3109 = 128'b11000111111011100010101111011000100110000100010100110101111001100000111101110000111100010101100000101100010011011101100100100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3109[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3109, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110011011000011010010101110000001010001101110101000111100111011001100100101010111110001101010011101010000010001111100010001110; 
out3110 = 128'b01010010110111000011101101111000100110011001001000111000001111100101000101101110100100100001000010000001010001110111101111101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3110[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3110, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110011110011000001100100100011101111110010111111000001001111011100010110100100100110101010111101011111000111001010111000011011; 
out3111 = 128'b01101110011100000101001010010010001010110010000101001010111010001100010011001011101100100010111110010000101101001100110111010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3111[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3111, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001100111001111110100111100001101001010010001110101110000000101000110110100000110000001001011001001101001100101110000101100; 
out3112 = 128'b11010001001001111000000101100001111000111000111000000011000101100110110110010101010010010010111111111111000100001010010000001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3112[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3112, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111101011001010111000010000111010010011101000001010111011100100010011011101100111110110100010001001111000100001111000111111100; 
out3113 = 128'b11110110011110000000001101000111110111101010001000001101100110101010001001011101110111011001101111110010011000000000100111110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3113[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3113, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101011010001001010010011011000110101111101001000111000111101011001111011010011011111111011110011010010101010011101100000001; 
out3114 = 128'b00001010110011001000101000011011010111100000000010100111101110110111001001100110010001110111111100111011011010010001100001001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3114[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3114, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011010101100100111001110110000111110010100000001100111111011110111000111000101110000100001101111101111101100100101000100100; 
out3115 = 128'b00101000000000000011011110001110000010001001011001000011000101101011000110100000111011111101100000001100111011010111101000011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3115[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3115, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101011100111100110000111000101100110100110001011110101110011011010001011000010100111101100011001011011110100001111001011100; 
out3116 = 128'b10110101111011110000001001010011100101010011010101001000011100101000110001111010000100111001110000010111011000110000110001010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3116[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3116, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000110101110000011110011000010001000111011001000100110010110011101110011011011100111101111010110110010110011010100111010101; 
out3117 = 128'b11111000101100000111101110100011100101110100101100011100111010110111011011101100010000011000110100101111101001011100111110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3117[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3117, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001011110111010111110010010001110101101001101001001010010010000001001111001000111010101010110111101011001101110100000011000000; 
out3118 = 128'b10001001101110011101111001100001000101010101011110000100010000000000000101010011101010100111100100000010100100010100010010010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3118[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3118, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101110010000100110100011011011101011101010100101001011010101100110001100110001110111100001000010101111111110111011010001110; 
out3119 = 128'b01111010110110011110110101000101110000000100010110101010101101111011010101011100111011011001110010111011111100011100011110010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3119[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3119, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110001001110000110110111101010000011011011101011010110100010100101100111000111010001000100101100000000100011010111101101100; 
out3120 = 128'b11110111000101001001100000010000110111110011010001011101111110101111100011010010000011011000000110110011011111011111101010110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3120[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3120, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010001010000111101101010000011011011000000001001000101111011101101001001110101011000100111001101111100100010110011111010101; 
out3121 = 128'b11100011101111101011000010001001001001010100010001001110111011100010101000000100001011101001001010010100000100010101100011110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3121[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3121, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001001110011100000101011000101001110111100000000000111101000100000101000010101110100011000011010011001011010110101010100001; 
out3122 = 128'b11001011010110110101010110010010000011001101000111101001011010110011001110111101000100100111001010101111110111110011010110101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3122[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3122, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000101001111000001111010110011110011001011111111101110100010011000100101101100010010011000100010101101010000110000110011110; 
out3123 = 128'b11100100101110001101101011011110111001011001101100010001011011100101101110110011011011111101100111101111000001011001001010000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3123[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3123, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000101001001011000110101111001010001101010010000001010010101100111110101110111011110101101000000110001001011010000101001101110; 
out3124 = 128'b01100111110000010011011010000010111101000001011010000000011001100001011001010010001110111111011101111011100001001100011101101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3124[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3124, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010011101101001001010011101000110100011000001011111101101100110000000101010000111010110011011011001111101000011001111010110; 
out3125 = 128'b00110010010100100011000101000111011011001111101000011001001100010110001111010000001011110111100000110101101001111110110001110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3125[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3125, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010100001110100101100010000011010110001100111110000100111110011111100000001001100001100010111110110101001000001011110100011; 
out3126 = 128'b11100011111011000010010100000011101000100101110110010101011000100110001011011110100111011101010101001011100010100101110101000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3126[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3126, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010100100010011001010000000101111000111110010111001100001110010011110001101110000000110101101100001110100111010000110000000; 
out3127 = 128'b01111111111000100011101111110001111001011110011101000101011000110110101110100110010101010001111100100110110111010100110001101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3127[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3127, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110110100110011111000001110110101000001011111110011100100001011000011100100110110110010101100000011100010100100000100000101; 
out3128 = 128'b01101110010011011100001001010110010010100010010010110100100011110100010111110000000001000101110000001111110101001010010000011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3128[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3128, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010011011011100110011110101111100111010000111010101001111011010101001111001000100101110000101011111100101011000111000100001; 
out3129 = 128'b11111101110100001010011110001000010011110000100010111010001011011011011001011001011111110111110101000001000000001000001000100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3129[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3129, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001000111101110001011011000001100011011111100010110011011100101100100011101001000110001100000101111011100000001100000101111; 
out3130 = 128'b00010010011111011110001011111110010010101110011101011011110111110000001110111011101010101101000110000010110000000011011110010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3130[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3130, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001110000110011111111101111111111011111100110011101100101110010110000101110011110100001011111110111011011000101100000010110; 
out3131 = 128'b00111111110110010011110101010010011111110101000000011000000010000100001000010111011010110100000001110110100101101011110011111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3131[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3131, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100000110010111000101110001011111001011001001111001100011111101010110110111101010000011000010100111000101111011111101111111; 
out3132 = 128'b01110001110011110101011000010110110000100010110101001110000001101110011011101010110001001010110010100111010101100100000100111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3132[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3132, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011001111101100100001110100000011010111010001100101011100110010101000010111101000110011110000000111000000001010000111101101; 
out3133 = 128'b10101101110101110110011010100101100111010101111101000011000100001001010001111010111000100111111000000001111111001111010010000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3133[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3133, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110111101111101101100000001111100011110110001000010110000101011010110101111110110110101110100010100010101011100010010011110; 
out3134 = 128'b00110111011011000111001110011010000100010111011101001100110100011110110110000001101100001100010110101001111111100000000010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3134[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3134, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111111111101101000010011100001010110011110100111010111111110100001000010001001001000101000000100100110111000111100001100001; 
out3135 = 128'b11010010110111010010101110010011011101110010010100010110010110001001101111111101010110101010000110000000001001100100001101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3135[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3135, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010001000111010100111111100101010101110011000001001000011110011001111100000101110111111100101100000001111100000011100100101; 
out3136 = 128'b10111111110010001111001010001001001100001011001111101011001111010000110111001000111101100010001111001111110001111010110100000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3136[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3136, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001010001010010010011001111011101010110000110000010001101011100100100010010100100100000100011010001010010111111010000010101; 
out3137 = 128'b11110100001000010010011001010100001000001001001111010100001100001110001101010111001110101001111111011000110011000001000000110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3137[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3137, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100000011110011000001110011110110110111000011011101110000111001010101001111100010101010101001100011000001100111000111000110; 
out3138 = 128'b11100110010110000011000110001110010101110000100011110111101101101010101101011010110010110100110101110000011011001010110110010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3138[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3138, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001111101101111101010110010100010111111011101111010010010001101010110000100101001001101011001101110000111000100101101011100; 
out3139 = 128'b10011011101010001111010001001110011001110101001011001010011110010000100100011101010101101111110101101101111000100000011110101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3139[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3139, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101001010101001110000101001101100010110101100011110001010101101000001011100001001010100001111010110000110001100011110000100; 
out3140 = 128'b10110011000110010000110010110011000110000110101010111110000010101101000000101000100000101000110000001010000000000101101001100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3140[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3140, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010010010110000010111101000101010100110111000110001101110000110010111000001110011000101111111010001010101101010100011001001; 
out3141 = 128'b10110111011111011100011111001110000100001100001001010111111111101010001011000110000010110111011010011011000000110110000011110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3141[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3141, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000101110111100001100110011100000101111001011111001111100101001000111101100110111110111111010000001011111110000010110100011110; 
out3142 = 128'b10010100110000011111110101111101000111110101101101101000101100100011111111000110011010110000010000111101101001100001111101101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3142[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3142, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001101010110011110010110101011101110100000111110101110000111000000111100110001011001000100010001101010110001011101010010010; 
out3143 = 128'b11111011001011111100011100001100001111001111010010101110110100100001010101001111101010000110111000100101111110101010101111001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3143[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3143, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110101011101111010111101011010001000000101011010000000010101111110101011000000111110011111011110010101000000110101011101011; 
out3144 = 128'b10101101100110011101110101010100111001010110110100000101110100110101101001010000101110000111001011111111000001001111100100100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3144[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3144, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011101001011011010001110011110111001011000010001011000001010001111001110011010110001011100010010100100011001010111101010010; 
out3145 = 128'b11111101101001110000110000011000010010111011001100000000111100011101001001010100011011000000111010000010011110010111110110000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3145[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3145, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000011000000110101100000110011101001000111010111101110011100101101000100000000000010000100000110010000010101001110110010010; 
out3146 = 128'b11100100011111111010111010111011011011001001110100110100111011100101000101111001111110010011101011101010110011010101111001110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3146[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3146, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101100001011010001101010100100011110110010111010001000010100110110011101101011111101110101010000010111111000010000011011010; 
out3147 = 128'b01101011001010010101111010010110000001011010000101011011000001111100000000011111011111101001010111011110011101101100111000101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3147[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3147, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011111000110011011111001011001001001111000010111000111001110011010110011100101010110100000111000010011010100010100000110110110; 
out3148 = 128'b11100101010100011100100000111001001100011110110100100001001011011101010100110111010100011101001010110010010110100000110011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3148[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3148, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110101110001111100110000010101110111010001010000011011110011000011000000011101101111101010011000101011001001000100011011011; 
out3149 = 128'b01000100111101101010101010011101111011110011110111000010011101000110000110010011100100011011001111001000100111111100101100001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3149[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3149, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000111111100000011001111100000100110010001111010001000001110001010101001100001100100011110000100100000001100111101110011111000; 
out3150 = 128'b00101011100010001001111011001011101001100000110100010111000101011001101100110010110011011000010100101011101000010101101111100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3150[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3150, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101100010100000000101001100110001100100100101000111101000011010001011010010011100110101001011100011010011000110011000011101; 
out3151 = 128'b10000001111000110110010010011011110100101110001111000011110001001101111000001001011000011001100011001010110111111001001110001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3151[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3151, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100001000101011100110101101000000110100000110100000011111101000100010101110001110010010110010001110100100101000110001110010; 
out3152 = 128'b11100101001110001010000101111011001111010000000010011000000010001010110110101101001110010001000101000101001010101010101101010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3152[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3152, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000010001101110011111100001110001001011101100111111011010010000110011111000101011001110101000001001001110110100100001101100; 
out3153 = 128'b10101010010001101000001010000100011111011010100011100100101011101111011101000111100100110111001101011000100011000011110000011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3153[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3153, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111010111100111110011110000011100110010101010101011011010010111000010000000000011001111111000001101110010000010011110010011; 
out3154 = 128'b10011001100001111001111011001101010011001111001111011111010110000000001101110011111000000100100001100110111010111100101011010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3154[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3154, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001010010010110100001011010000010110101000100001100001110000101100001100011110101001010100000010001000101000001101111101101; 
out3155 = 128'b10000010100001011000100110110110110011101111001011000000101011101111110011111110100101110011110001110001101000101111100010010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3155[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3155, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101011110001101000011100100110101110100111000110111100001011010000001010000001000111001001110000101000110011111000011000110; 
out3156 = 128'b01110110110101001001111100001010000100111010111001101011000101111110010111011101100000000100110011110001000100110111001110000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3156[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3156, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100010011001100000111110110100101110110101110000100101000011100100100001100011100000011110010100000010111101110111101000100; 
out3157 = 128'b00000100111110011010110001000001111001010010010001101000011111101100100111010101111011110100100011011100001001011100000111011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3157[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3157, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001111111010110001101100101010001010001100101010110001000001011011101001110100101100011010101111100000011111101010000110110; 
out3158 = 128'b10101101100111010110001110001111010100111100011010111110111000111001111100100010001001100101110010001011001101111110101001001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3158[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3158, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010010001100101101000111110011011101010001011011011010000011001101111010010001110011111001011010110111100111100010111110110; 
out3159 = 128'b11000100011100110101001000010110000000101011100000111000011110110110110101110010000110111000111000111101110110011011000011101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3159[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3159, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101100001111011001100001010100000010000001110100110111011000000111011001001001111001010101111000010110010101111011111010001; 
out3160 = 128'b01110111011101001110111110111000001101100111011111111011100100000000011111001100100011101110111011101011100001101110010000111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3160[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3160, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010110110100010011001110010100110110001110101110000011110110011010000100010111101011101011101001110001010000111111001110101011; 
out3161 = 128'b11011100010100000110011010001011001111110000110011011110011100010001100110010000000010100000000111101011001110110110000111011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3161[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3161, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111101100000110110100111100100000100100001100001100101010111101101001101100010111000110111100111010011100001001001010000110; 
out3162 = 128'b11111001110110011111100010100101110010000111000011010000100010010011001110100000101010010000111101100110000110101110111001000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3162[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3162, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100011100000001111000100101100110110010000010001100111011000110001000101101011001101000000110101010001111011000001001111001; 
out3163 = 128'b00111101010101101001101000001101001010111001010011001101010010011100010000010110100000001101110001110011110010111010110100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3163[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3163, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011011011101111001001111000000110000011101001001001111001110110110101011011111000101100101001000011110101001100111111101110; 
out3164 = 128'b01111110011010110101000100101111100100011110001110111000101010011001011000101100011000100100010011110101111110101110011000010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3164[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3164, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111101110011101000101010100101001010011110110110111110101100010100010111101010100101001010011000110001011100001011010110111; 
out3165 = 128'b01001010011001101000111110111110100111011001101101010010011110110101011100111101011111111111001100000100010011110100010111010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3165[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3165, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101100110101100011110111000001100001000011010101011100001010011100100101101001000111010010100000111001110110000101101111010; 
out3166 = 128'b01111010100101111001101101000000100000111100110101101011001101001100110010001110111111101111101011000100010010001011100111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3166[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3166, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100001011100001000100110101000110011100000100011111011010111011101011010100110001111110000001101011101011111011001101101101; 
out3167 = 128'b01110111001011101101000011001100110100000000111000010110001111001000100011110110001100001011010000111101110011001110010110010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3167[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3167, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100101110111011101100010010100011111100010101000100101100010100000110100110111001000001111111000000010001011110101110111111; 
out3168 = 128'b00010010000101100000110011010101110011111111100000000100101100010001100001110111010110101111001110010000111101100111101010010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3168[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3168, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100111001111000101011100010111011010010101111010110101101001010011101110000000010110010111011110100110101100000010111100110; 
out3169 = 128'b00010110001011111110011010111000100100011100111001100100101001100010110101000111011000101111111101111001100010001100011011010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3169[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3169, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000000010101100100001110010001000010010110111111100001011100011011011110111011000101110001110111010000001110001110011011000101; 
out3170 = 128'b01101011101101101110011110110100101000100010101111000010000111100101010100110101110100101100010010110101001010111101110000011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3170[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3170, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110011101110010011100110001011101001111101010000110100011000111111100011000111110101101011100111011111010101111010001110011; 
out3171 = 128'b01000011110000100100010100101000010000100011001001001100000110110000111000101011111000100010010000111110110101111101101101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3171[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3171, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011110101011000010000000101110111110011110101001110100010100100001111101110010011011011100001011011111100000111101001010100; 
out3172 = 128'b10011011111110100111100010100110000000010100101111101001100110011010111100011001111011100100000001001010100010110010110010011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3172[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3172, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111010000111010001010011110001001000011101101011000100111100001011110001100111110010000100101101011011011000001110100001010; 
out3173 = 128'b10000100101110011110011000110110101000110000100111000000011000010000010001111111101101001011111010001001100111001010101001110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3173[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3173, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000011011011000110001100101110011001100101001001100100010001010100110001111100101110101110110100110011111111110110010001100; 
out3174 = 128'b11001101100011001001010101111000001000100110011110001101111110111010101011011101000111000000010100011011010111001010100010110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3174[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3174, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001100110111010000111011001011111110011101110100011011010110000010100100011000111110100000000100011010101111111000101010100; 
out3175 = 128'b10001100000000101001000100011101000000110111010011001000011110111101001000000110010010101010110001000111111111100101111101010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3175[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3175, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111100100100110011101111110010101000000101010000010101110001100111100110011010000000000000101101010101111101000100100110010; 
out3176 = 128'b00100101101001010001011000010101011111100001100000001101101000011110010001010111110000100101110101101011010000110011100101111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3176[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3176, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101011100001001101000101111000100000010011011101000100110110011011000001100001011110011110111110011100101000110101110100011; 
out3177 = 128'b00000111101011111010000111101000111110110111100111100011100011010100111010011101001000000011001110110111111011001001001100100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3177[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3177, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011101010111011010111110001101101101011100010100000110110000001101100000111101010011000110100101000100010010111101001001111; 
out3178 = 128'b10111101011101111101011101010001000111011101010000101111000101011000111011011011011110110010001010010011100011101110000011001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3178[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3178, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110110101110111001110100110111100010110000001110000100000001001100010010100010011011101100010111111111100010001100100110010; 
out3179 = 128'b10110010001001011011100000010011110000101000011010001010001111110011110011011101001101010111101111000011110011101011001011110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3179[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3179, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011011010101111000100011111100100110111010001100100101100101100110001111111001100101101111101000101111100110110010000111000; 
out3180 = 128'b00100110001101110110011010000011100011110101110100101111100111111001011000100000111100000001100101011001001110000010000110000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3180[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3180, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110000111101000100100000010010101111110000101000111010100111110011111111111101010001100011101011011011001010010001001100111000; 
out3181 = 128'b00010110000111001011111010001000010110011111001001100111001100010000110010010000111011011000011000101011010010101100100010100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3181[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3181, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001100101111001000111110011001011011100001110011000100101001111101111011011011011100111010100101001010100110110100101111101101; 
out3182 = 128'b10100111100110111011011000101010100001111110000001111001110011101110101000011100111001011100101001001111000010110100110011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3182[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3182, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001101011001101000100111011101110100110000011000100011010101110101110101100000001010100111001000000000111100111011100110100; 
out3183 = 128'b11100010110000011100110001111110010010100010111101010100110011110001010111001110010111000101001111100010100100011010010001001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3183[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3183, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010101100011011011011110001010100101001110100101100000111101101000001010100000111011101100110100000110101011010000001100000; 
out3184 = 128'b00000010000010101000110011010001100011001001100100000100001011001101011010111110001011110000011001111011000010101111010101101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3184[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3184, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100010010101001000000110000101111000101000101100001101111011001100101101010110011000101000001110110101101101010110000001010; 
out3185 = 128'b01000111000000110101110010110100111011111000111110111111001100011000100100111001011001111111001011111100010100111011110110001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3185[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3185, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111010111100111011001110111001111111011011011000100001011010011000000110100011001000011110001010100010011110111101110001001; 
out3186 = 128'b11001110111101110010101001101000101110100011110001011011010001000000000000110011001000100110110010010010101100100010100110010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3186[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3186, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110011111000001100011000110011100110000001100001100010000101110011001101110100001110100101100101001010011101010001011011110; 
out3187 = 128'b11000001011000001000001000001110101010000001110011101110111101001110111011000000101000000000001111011001101100110001110011010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3187[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3187, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011010100000100000101010111010001001111010000101110110100001100111010101010101111011000001111000010001100011111101001000110000; 
out3188 = 128'b11111101001001111000111111111111010101010101011011101011000011110111100010010001101001101000010001001000001110101011110111100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3188[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3188, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001110111001100010111000110101011010101001110011010101101010111000001001110100010001110000100110111000110000011001011100110; 
out3189 = 128'b10100010011010000001011111110011100010010010101100010000011011110010100010110111101111011100000000011011011101111000101110000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3189[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3189, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000111001111111010001111001000100011100101111000100010101110101111100100010001000100011101100101110000111110110101100101100; 
out3190 = 128'b10000110101001000000110110110001010110000100101011001111101110001100100110111101000001111111111010111111010010011011111011101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3190[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3190, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110100001101010010001000001110101100000011101100000110000001101101000101110001111001010011000110010101100001111101011110001; 
out3191 = 128'b11101001110000011110100101100110001111100010000010101111010001010111111001000111101001111111101001000101101011111110110110110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3191[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3191, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010000110101010111110110001010101100100100111110101001000000001100100001100111000100110111010111010011101011100111000000010; 
out3192 = 128'b11110001101011001101111111001011100110101001011001111001011001101111111101010011001101011110010110110110011001011010100010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3192[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3192, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010001100011100000111011000100010110000111110100100000100101100101000010101101101001111100000111100111010111100011001000111101; 
out3193 = 128'b01000101101011001100000111110011001111110000001011101000111001011110000101101101011111000001000011100001111100001011111000110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3193[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3193, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100110101011010011110101000111111101100101011101000010110100100100100001111011101010010111111011100011011110000010010111010; 
out3194 = 128'b00000000001110111011001100100101011111001100010101101001111010000011000100100011011111101101000001111100111110101011001110001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3194[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3194, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011100101111100101111011001011101110010111000000101010011000110111001101010001110010100110100011101011101010010011001111101; 
out3195 = 128'b01011000100000100111001011100000100111001001100110010010001100101111111101101111010110100000111101010101111010101010011000011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3195[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3195, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111111000000100011100111000000001010111000000110111000011000010101100111100101000010000100000110110010000001010011001011100; 
out3196 = 128'b10010010110011101110110101001110101100000000010000111000010001000000011111110000110110001101000011100100000101111010011001011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3196[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3196, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101101101111111001000000001001110101110010001011011010011001111000000000000111011101101010110101001001110000010111111000110; 
out3197 = 128'b01010101111010101101010001011111010101000100010011100100000001010111111110001001101000010011001010011011110001001110110100000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3197[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3197, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011000110000010010011011011010001101011010111111001001011100011011100011010011000100111110101110011100001001011011100100001011; 
out3198 = 128'b01011111111101100001010000001001001111001011000011101011110110111101110010100110010000101001011111111111010000111000101010000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3198[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3198, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001101010110010011000000001001101100011001110001010101101000101010001001100111000100110111101100010110001010101111001000001101; 
out3199 = 128'b10011110010110000011101110111110101000110000010100010110100011001001100110010110101000100100011001011010101000000100101100110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3199[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3199, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101011000101011110100000011011000110011101000100010101010110010010000101101100110001000100100100111101011101110111000000111101; 
out3200 = 128'b01011111111010000100000010111100100000100100100010010001010101000010010011101111100010110101111011101101010000111110001111000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3200[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3200, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110011010000101010010101101111001111111100110011000110010001001110001001111001011100000000100001110010010000011010001111110; 
out3201 = 128'b00100100011111001110101100101100101101000010111011000101111001000000101110110011011101110111111100100000100101110101001100001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3201[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3201, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100110001100010010001000001010111111001001001010101110100010101000010110010101001100010101011101010001101001000111010001000; 
out3202 = 128'b11011000001010011101100110110100001010110110000101001011101110100000010011111100100101011000011111110100011111100110101110100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3202[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3202, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100100011111101000110011111101000000100101001101001100000110000111100110001110000000000100110011101011101101110010100011110; 
out3203 = 128'b11010100110011010101110000001001101100011011110001010001011000010111101011100011100110011100001101001001100111111001000001110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3203[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3203, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001110000010000110100101000111011101101110100000010001101011101001111011100101011110111111110011110011001110100100101011111010; 
out3204 = 128'b10111101001000100101010001001101100001101111101101101100010000100101101101110000001100001101111010011011100100101001100111000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3204[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3204, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110111000111001000010111111100011000001000111100100111101001001011110011011100100010010100110101011000001011000100101111100; 
out3205 = 128'b11101000100101100011001000010111101010101011110101000000101000101101001000010001101101001110110101001011100000111101000100110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3205[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3205, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001011011110101100010110100000101110000110000111010101111000111010111111001001110100001100110000111011001001101011100010111; 
out3206 = 128'b10000001001111100100000110001000010001100011011100101111001110000011001000110010001001101111101111011100000011010000110010011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3206[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3206, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100001100110001010101110111000100111001011011010110011011110001010110000011000011000110010001010100011111000011110111001011; 
out3207 = 128'b00111011011100100010000010011110101010100100011110000000010101101100010001011111011111100010011111101110001110110000010110110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3207[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3207, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010010011011000011110011111000110011011000000000100010011000000110000111010000010100101100110110001100100110000101010000101001; 
out3208 = 128'b11100100111111111110010101011100001110111001011110000101111000001101100011000010000001001111001101101111111100010010000010111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3208[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3208, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010001010001100000110001111100111111000111011100110011010100000010111011001111111110101111011111101011001101111010010010010; 
out3209 = 128'b00111101010010000001101001100110010001011000001011000110000101011111111100101000101101000101100011100111011101001001001110111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3209[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3209, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010101111001110110100111010101010000011011011110001000111010000110001000011011110000000011000000011101001111111111100101001; 
out3210 = 128'b11001000010001010010100001001010001011101000101110100111001100110000010110101011010000100110001111110001010010000010110011001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3210[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3210, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110001011101111001111001001011110011111101010001110100010001101011100000100001111110110000101000111100100001100001111110111; 
out3211 = 128'b00000110110100010011100110010010101001110100100001100000101000100001101011001111110010100111000000100010010111101000011100100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3211[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3211, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001001001011000001010011001010010000010100010111111011100011001100011011011111111101010010110000110110110001001000010101011; 
out3212 = 128'b10101011011110011000001010010011100110100001111011110110100000001110010001011110111011101101100101011100110010110010010000100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3212[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3212, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101100111010100111000100111001101000001000000101101111010001001011011001100101010010101010111101011001011010101000111101110; 
out3213 = 128'b10001110000110000100010000000101011111110001000111111100111001101010110001000010010110110011100001000111100000111101010011100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3213[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3213, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000100101111100000101100001001000101111110100001000100101110011111111000001100110000101100111111011110110111101000101110100000; 
out3214 = 128'b11110101101110001100100011010001101000001100000000111011010110111001101111110001111011010101100010111010100101001010011000010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3214[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3214, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101001110000111100011011110011011100110101000011011110011000010110100101101100100101101001111000000010000111000100110010111; 
out3215 = 128'b10010010111001000000111010110110110101100111101110010000011000100101111001000011100000110010110111000010101101011000101001111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3215[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3215, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000001001111101011111011010001101111011000110001000000100101110110000000010000010001011000010000101000101011100111110111100; 
out3216 = 128'b11100000100111000000110011111010101011101000110100100111011011101110100111011110001110010001101001100001111011001011111100111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3216[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3216, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100000011001111111111100000101100110101100101100011100010110001010101001010100010001000110000100001111100100110101001000011; 
out3217 = 128'b11001111110101011110000111010011100110110101110100010101010101001000001110000111011011111001111100010110000001101000011101100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3217[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3217, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001100100110101010100010111000111001011101001001011110101011011010111000010010011100111000100101001100100100101001001000101; 
out3218 = 128'b00000101011000110100010100100010001111111000100001011001101011000010001000100100010011110100000101110110101101101101000100000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3218[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3218, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101111001101000001000111001010000110100100111100010011110110010101010110011111100100111101000001010010000111100100111000000; 
out3219 = 128'b10111100011111101101010011101011111111010011000011011010011010000100001010110001001001011010110111110110011110010111111011011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3219[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3219, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101100111111011011001011110011101000000100010011011000010001101001101000101110110100101001001101010100001010101000001110111; 
out3220 = 128'b00111001010000011100111010101011011110001001111111111000101101100010101010010101001101010011110111001011100010111001111000001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3220[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3220, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101010111110110000111100010110010011100110110100010101101011000001101000001010000000000001100001101100110000110110101001111; 
out3221 = 128'b11011111000100011000111110000000110000111000111100110100101001000011001001001001101111001110000001101001000100010110001110111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3221[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3221, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111100011000101011110100101010011000101110110010111010110100100011001011011010010010101110011000000011100110111100101110101; 
out3222 = 128'b01110011110100010100111111100100100111101010100111101001010000001111010010111010100000000100110101110110000001110110001100000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3222[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3222, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100100010011011010010101100010000100100111100100001001100001011001010010100001100011001100001101110110001011100001000000110; 
out3223 = 128'b01101110010001001001011001110101111011010100110100100110001110110011000011011001111001101110010110110101110011101001101001111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3223[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3223, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110001001100101010111011111101001111011000100001101101011010100111000011001001011000001011110110010110000110110000100011110; 
out3224 = 128'b00010100111110101001110101001011100000101011110101101000001100001100000010010010110000100011110100110100000100001011010010101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3224[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3224, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010001111000101011110111111011101110000111010101010100001000000110000100110101011111010001010111011100000010110001100011001; 
out3225 = 128'b10111001001100011011000010100001101011001110011000111110000001000001010100101100110110000011100001010111010000101110110010010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3225[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3225, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110100010010001111111101111010001110110001110001001110100001001110111001110011100001101100100001111111011110001101000011000; 
out3226 = 128'b01010001000110111100100001111101011111101111110100101001111100110100011011110011110010001011101010111010000101110111110010011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3226[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3226, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111100001110110011111111001110100000100010000001101100111011000110111100101101100001011000010000010000100000000101011000011; 
out3227 = 128'b10010000101000001111101111100011001110101101010111010100100111110101110001100110011000111111110000100110011110010100110110101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3227[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3227, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000101101001000111110011101010011100011101000101110110101011110011001111000001001111011100100011001100100000100001010100000; 
out3228 = 128'b10001110011111101101101110000000011111110001101100011111111100101100011011011110011011110100111100010010111110111111010001011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3228[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3228, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110110000011011111110110100001100010011000101101001001111001100100010001010110001110000111110010101011111001000001010001001; 
out3229 = 128'b10110001010100011011110000100010010010010001001100000010110010101001111011100011011111010001001010011000010010110110001000001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3229[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3229, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001110101010001101011001100000101110100110001101011101111111011010101100000101111101001010111110010011100101101110001111110; 
out3230 = 128'b00001111010101001000100001010100110001010001110100110101100011101111101110100101001110100010011101111000011011000110000010000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3230[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3230, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101000010001011010111010100011001101111100010011111011100100100111111011011110010010000000100010011100011110100000100110001; 
out3231 = 128'b01100011001110000010000100011000110110100100101111110100001111111001111110010111110010010000000010110000001110010110001001001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3231[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3231, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111010011101010010110000010101100100000110100010010001100100101011101001101001100010111101001100111110011000111110011110111; 
out3232 = 128'b01001000100010101110110100110001111100100011000111111011111001110010100100010100010001010100001000111110000110110001001110000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3232[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3232, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001001100100000000110110110000000001101101001111101001101000111101111101110110010100010010100100101111000110011001010000010; 
out3233 = 128'b01100000010101110100011100011100010001011101101001001011101010001110110000001110000000011100100110010100101001011011010110100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3233[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3233, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011000101001010101101110011111010001011000100001010101000000000011111111111110010001100110000000011001100000001111100100111; 
out3234 = 128'b00111110010111010110010000101010010110000001011111010011010101110011001001000101011100010010010101110110110100111001011101111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3234[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3234, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001001110001011111010000100101110111010111101010101000011110111000010110111001001110111110100010110101001101100100111001001; 
out3235 = 128'b10111000111000000110001110111010000000101011010101111010110111000000001110001110111100011000010100110101101110111011110011110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3235[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3235, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111110110000000001011111010000101110100010010110011100011111011100001000000010010111111100010110010100110101001100000111000; 
out3236 = 128'b01111000000011000101110011011111011000010111001111001110110100000000011111000101100000001010001000001000111110001000001001010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3236[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3236, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100101101011111101001100100011111011011001110111001010000110001000010010101011101111000001010101001000011010100001011001000; 
out3237 = 128'b01111010000001001001011010010011110001110011110011010001101000001001111011000000101010111011000110000001100111010110010010010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3237[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3237, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100010100110101101011010000111011000100100100101110101001111111101101101010000000011111001110111001010000111110100000001100; 
out3238 = 128'b10011110110110000100101100000110110101111001001010111100001101010111011001100000111101101101001011110001101110010001101100110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3238[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3238, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010011101111001111110101101010101001010111011011100010101101001001001001000011000000000110000010010001011010101010000001001; 
out3239 = 128'b01111010000111000011011001010011101011010010101000010111001101001011101011101001001110000011111000110101001000001001001011111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3239[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3239, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010111010001011000001111001011110010100100001010010010001000000110010111000111011101010000010101101110011111111110010110101; 
out3240 = 128'b00111011001000111100011100011101111000010100001110000000100101111111110011011011001010001100110010001101000111011001010001101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3240[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3240, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110001110101101111110011011101011101011010111000000101010010010101011110100001011000010000000110001110000010011100111101001; 
out3241 = 128'b11101110110000110011100100101101100100001011100001110100111000110010101010101111011111011000110011010010101110001101000111000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3241[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3241, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110110011101001000111001011101100001001011011010110000111000000111001010111110011011101101000101011010101101001011011110001; 
out3242 = 128'b01001111100110100000110010001000001100001111011001011100110010101010000110101110100101110110100111111100010001100000001010010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3242[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3242, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100111011011000000110101010011000001110011010101100011110100000110111110011100100100110111011110011010010000010100101001000; 
out3243 = 128'b01100011100001101000100101001101111011100110101000011011100010111000001111110101100000001100100000001100011010011100011001000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3243[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3243, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100011010000000000100010010110100111111011100111001100011111010001110010011111010000000011001110101100010001100000011000100; 
out3244 = 128'b00010000001111100011000001101111110000101101100101010000001100101000001011101110001011111000101100000010110011101101010011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3244[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3244, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110011000111001000110000111110000101000111111000110011100111000001011100010101011001001011110000101000111001011101001010001; 
out3245 = 128'b01011110010111010011100110110010011010110011011110000010101001010010101010010010000010101100011010100100111001100111011001101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3245[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3245, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000001101110000111110000000110011000011100110010110110010000111110010110000100111011011000111111010011100001101000010000110; 
out3246 = 128'b00001010100111011101000111001101111101000000010101000001100110000100110101010010110110010010100110010001001111000101110000110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3246[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3246, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111101110011011010111111001101001011001101010010010010101011111000000101010111111110100000001011101001100110010000000011100; 
out3247 = 128'b01001011111100010110111011010010010001010111111010010000011010110001001010010011101011101001111000110000101110001111010111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3247[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3247, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101111011000011000001101101110111010101101010010001010011100011101010110110010001111010011111110000111110101110100111011010; 
out3248 = 128'b11001101101101111011001001001100111100011100001100011101000110111001010100110011100000100001001101000101011110010001110000100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3248[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3248, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101111111100010100011000000001110000110011010101111111010000010000010000111011001111000101100000111100010111110000100110010; 
out3249 = 128'b00100010100111110000101101111100110110010001000101000001000110000110101100110010010101000001100001000011000100101111000010100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3249[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3249, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010111110010110011110011010100001101000111010111001001111111011000010010101010001100010100110011001000111110001001110011011; 
out3250 = 128'b11110101011010001001100000000100001100000101000111000110111001010111011110011001010101001111011110101000111101101100101111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3250[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3250, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100111001110111101110101110000111111000001000011011100110111111001101000010011011101001111001010111001110010111000001100100; 
out3251 = 128'b00011000010011001011110101101101000011100110000001000000011101101010001010000110001001101011000011000011010110010001001110001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3251[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3251, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011001010100100111111001111110100101111100111111011010011100011100100001111101101001101111000100000001001101010110011010110110; 
out3252 = 128'b01001011011000111101110011000110010011100111111110100010010001110011100010111000111110100100010110011111011011001011110101010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3252[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3252, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011100000011111011011111011100011100111110101101010111010010111111010000110100011010100001100000101110000111000111010101100; 
out3253 = 128'b01011111101011010001101101101010111111001001101111110010101101010011010101011110000100100101011001010111001010111011011001011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3253[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3253, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111111111011110101110001101010111110110100111000110111111001011110011011010101101000100111110110110101000111110011010001111; 
out3254 = 128'b01100010100001011100000101100010100010000000000010001110001100101000111111011110000010000010001001010011011101110011101111010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3254[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3254, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100010000110100110000000000101001011000111000011011111111110110000101100101011011100101001110101101001000110011101101110011; 
out3255 = 128'b10100111101110000111110101111101011010111110101101011110101100110101011100111110101100001011001100011000010101010100111101110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3255[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3255, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001100011110110100000001011110011110111010110101110100101010011110011001010110100010010101110001100000101010011100010101110; 
out3256 = 128'b01000000001100111101000100110011111100111010010101100011100101110101010101010110011011101101010001011011111110001110000100111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3256[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3256, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101001001111001110111000001000100101001101111000000111100011000110010101111110011111111001010001111110011111100111001011111; 
out3257 = 128'b10000100110101011100101011001101001111110011001111101011111001111101111110101000010001010011011001010100110101011101001111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3257[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3257, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010000000010010010011001111001111001110111000100100000010011001000101100101011110011000100000110100100100100111010001100000111; 
out3258 = 128'b10100010100001100011001000011001111111110001011100011010101100110110001011101100010100100101110011011010000101011100101001001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3258[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3258, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010010010010010111001101111001011011100011110101011000111001011010100100100100011100111111010100111010011011011111101100011111; 
out3259 = 128'b00010110111010000100001101100111010010001000010101000101100011110011110001010011011110011000110011011111011111111000101100000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3259[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3259, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010110101111010110010000101001111011110111000010001011111011010011010110010100101101101111100000010000100000110100011000111; 
out3260 = 128'b00000101101000000001110101001111001100110100110000001100000000001011011010011011100111001100110000001000010100001101100110111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3260[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3260, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100100000101100101010011110111001010111011100100100010111000111100000011011110100100110011011110101111010010111001111101100; 
out3261 = 128'b10011000110110101111101101101110001000100111010101101010001001110010100011011100101001101010011010110111010110000011111001010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3261[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3261, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011100111110011000101010011101110111000110100100001111110111000001011100010000010111010110101110000110101100100110100101110100; 
out3262 = 128'b10111000101110001010010111010011010011101010110000101010000111101011011101000001011110110100101111001001011101010000010011001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3262[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3262, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111001110010000110011001001001011110111000010110011111000010001111001101001011011110101101110000010100011001011010000101010001; 
out3263 = 128'b00101111101001100100110100010100100100101110100100110000010010111000000000110000001110110111010011011011110110100010000000100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3263[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3263, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010010000100010111101010111011011100111000100111011001011011100010110110110111011000011010010011111111101001000111001001000111; 
out3264 = 128'b01110010111100011100110001010011011000110100000000101100110110011110111010101111101100000110111111100011100100000100001100101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3264[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3264, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110100100010110010111100111101110100010011110000100011110101001101111110010011111100011010011110110100100111101001011100001; 
out3265 = 128'b11000100000100110101100011011111111111001001101000000000011000111100110111100100000010010100001001001011010010101010011111110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3265[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3265, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001001011010000110100100101001101011110001101010011000100100100101110111000001111100011111001110111010110111110100001001010; 
out3266 = 128'b10101111000000000101000111001001001101100000100010001110001101110001000100000001111011011101010001010101101111011101000101000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3266[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3266, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000100000011010010111001011110011010000001100010110111100010010110111001000101000001001000001000111001101000001000110001101; 
out3267 = 128'b11111000010110100100100010100110111110111110011110011001010110101001101010111000100011010010111111101000101101001011101000010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3267[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3267, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001100000110100110101010100110001111110100101000001101010101010000100011011111111011101111111011100001011100100001110100011; 
out3268 = 128'b00110101010010001101100101001101001110110011111011001110001000000000001000010001111000111010110010111011100110110010101110101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3268[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3268, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100100110000110001110010100011011111101010001111001011101000001101100111100110100000110101111100101011110001001001011100101; 
out3269 = 128'b11110110011100110100100011010001110000111011000100010100001100100111110111110100011111011110000110100100110110111010111000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3269[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3269, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101011010111100001000010000101111010010001101010000010110001000110101100010010010110001111000110001111000011011101001110011; 
out3270 = 128'b00001011001101001101110010001011111101101010111111011010100011000000000010011011001000110000100110010000001000110000001111111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3270[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3270, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101000000111010111111110010000010111011001011100001110100001100010001101101111111011001001100100111010001011011101100101100; 
out3271 = 128'b01101101001100111100010000101010001010101110011111110000010101010011101101010001101011110011100011001100101011111100011001000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3271[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3271, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111101110010110110100110000101011101100100110010010010000001001100101001111100111100101101001011011010000110100110011110110; 
out3272 = 128'b00010011010111000010100111001000100111110110010010011100001000001101101111111011111100110010100001010100101011111101101100010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3272[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3272, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100101001111110100000011000000000010010001100111000011001010101000101011001100001010011111100110110001111100011001101100101; 
out3273 = 128'b01001101000000010001011010101110101111010011100000101101110001000010011000011101111011110010001111001010000000111101101010011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3273[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3273, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001110111010000101000011110110101110000011111010111101000011100111101001101101110000000000011111100110010011001001111001111; 
out3274 = 128'b00010110101100011111001110000100001101000000100001100100010111011110010100110100101010100100000010000111110010101101111100010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3274[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3274, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011011110000111110101001101010010101100110110111001010101111111111010001000110100010010101000111110110101010110100010001001; 
out3275 = 128'b10110011000001011010011101000001011101000010000011001011000111001011101110001001111011111001011011010000111100101000110010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3275[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3275, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011010110111000000110000101100011000000010011101000010110010001111110110101111111010001110101001011010110010110100000010101101; 
out3276 = 128'b11101111010101110011011101111100000001010001111110110010101110000001010110110011000001101100001011100110011000011010111011101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3276[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3276, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111010110110111001111101101000111101010000110001011001001111000111000111001101011100010111001000111010010010011010101010110; 
out3277 = 128'b10000000001100110101111010111010111011001001010101111100111101010000101110101011000101001010100011110010010011001000011011101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3277[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3277, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011100001001111111101110010110111100011001110010000111001101001100100001011110011000010101001010110101100000110111000100011; 
out3278 = 128'b01000101001110100011011110000110111101011011111111010100101011110110101010111010100111101011011110100101100101111001001000000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3278[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3278, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001010010100111000011010001111001110101000010010111111111000111010111111110010111010010101110011111001000110011110011001010; 
out3279 = 128'b00001111110000001111001010110001110110011011001110001100011110010001100101111001101110001110001110101011011001010000111000001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3279[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3279, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010010111000001111100011111111101010110110111011011010101001010001100001111111010101101111000111010010101101001001100011001011; 
out3280 = 128'b00111000100101101000010101011101011011000010010101010101010001011001100100100101101001011101110000001100011010000101100000101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3280[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3280, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111110001001011001000101011010100000011011001101101111110111101000001100101011010111101110101011100110110001110100111010011; 
out3281 = 128'b10110001101010111010101111010100000110011100110000000011100100101100011100011001001111011100110111010001101011011101110101001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3281[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3281, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110110010000111001101101011111001111100111011101010000011111110001011010011111001000010111010100110101000000010110100000111; 
out3282 = 128'b01000111111100010001000011101011110000011010001010010100100100010010001111110011001010100001101100100110000011010100101010111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3282[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3282, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000011110100110001011000100011111010001101001011000000100000100111000100011001101110100010110011101000101000001101110110000; 
out3283 = 128'b01100101111110001101001101011100101101001000000111101101111011011011001101011100000100100001001110110101010111100010001111100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3283[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3283, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010001100011011000110101010000001111001110100111001010010101001000100011001001010001010111010111011011011010111010100101000101; 
out3284 = 128'b00010010110111111001110111010111111011001001001011001011000000010000101100011000111010010010010100100011111000011010100111110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3284[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3284, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000010111100101011100011111000100000110010011101101110111010011100011011001110101110010000110000001000111010111101010111100; 
out3285 = 128'b11110100110010010011100111111100101011011100010000101111010101101011101000001101100111000000111100000111110110111110110000101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3285[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3285, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111000111101111011111001010100101000011001101011100000000001111100001001000001110000110111011110110110000001010100001000001; 
out3286 = 128'b10101100010111000110101101010001110001111110001011011010010111010001111001000110001100010111011101101110101110000011001000011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3286[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3286, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111000010100000111010100100010111010100010011010100011011100010000000110010001010101101001000111101100000001011000110101111; 
out3287 = 128'b10001000011111100111011010111011000011000111111101001110001000100111101110001000101111011110101110100110000110011000000110000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3287[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3287, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011111100111101110101110001100111110101011110110101010000101011101010111110111010010100110000011000110111010101000001011010; 
out3288 = 128'b10111111011101011000111010101111011111001011001010111010110001110011011110001011011101101111001101100001110011001110100000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3288[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3288, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111100111001011011011011001101111100000111110100110101110000011010110110010100101110101000000101011100000010001101111010001; 
out3289 = 128'b00100010101111111100111000000000110110010000000001110110110111010100101011110010110110001011011000001110101101010010010101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3289[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3289, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011101101010000111000110101101110110111100011100010001001111011010011010111110000110101110001111101111001010010011101111010; 
out3290 = 128'b00101100001110110001001010100010100010000000111110011011000111001101000101001111011101110010010010101010000111001010010100010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3290[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3290, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011110100111111111000101110001010010000000011100000101000010111011100011001000101001101111011101100000001010001111000001001; 
out3291 = 128'b01010110101100000010100110000000110110010000100001000110110101000001010011000000011010001011100001011000110010111001001111100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3291[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3291, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011111110101001001110111101110101001111001110110111011100111011110110110001000110000011001001001000010100100011101000100011100; 
out3292 = 128'b00110010101101110001101101011010001001001001000000100100010010110110011001111010100000011011011111000010111001001000000000001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3292[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3292, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001100111100001111000011011001010010010000111010111111100010001101000010010110100111111001010010111000101011010101011000111; 
out3293 = 128'b01100011011001011011001111011101000011101011111100101001101001011010111011101000001110110001110100011010010101111010000110101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3293[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3293, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101000001100101011000100110010010111011000101110001011000100010001010111011001000110001100101111010100010001100001111010100; 
out3294 = 128'b00010100000010101111101111101100110010001001011101001111101000100000011000011111001101010111100100000111010011001110000011110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3294[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3294, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111010000100001011100100011010110110000111110101110001100001100001010000100011010100111100001001101101110001100011000101001; 
out3295 = 128'b00111100111100100010101001000101000010101110011110101000010110110010010110100000001010111101100000100100101111101111010010001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3295[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3295, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001111111001100011010101000101110000011111010001100000111000001010000100101000111111100101100110101100000001101000110100010; 
out3296 = 128'b01101111110110101110110000000100111011000011001100100011110100011101001110011111100111101011000111001011001100110101101011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3296[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3296, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101110101110111001010111010100101100000101010100101100011100100010010001001011001001001111100000001011011101101001100110101; 
out3297 = 128'b01111001100110101111111101110011110000010111101101101001110100100001101000000110101000111100000010010101111110110010101011111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3297[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3297, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010010100000100100111111100010111111110000001010001101111110110001000011001000001111010110111101001111001001011001110000001110; 
out3298 = 128'b01100110110100000100001011001101001000100001101011011100001011000001001011100100011101000110001101111100111101100100011000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3298[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3298, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100111110101101110010011111001001000100110110010000001011001110011101101000011000011110110110000000110111011001010000000010; 
out3299 = 128'b11100110101001010110100100110101100111110010101110110111111011101001011110110011110101110000011110011100010110001011000000011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3299[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3299, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101001101111111100100010010101101011011000011111001111100011010011111000010000000111010011010101001110001011100111011010110; 
out3300 = 128'b01110110110010010111111000000110110010101100110000000011010100101110001000100001110101101010011111111001011101100011110111011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3300[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3300, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000010110011001011110111110101000101011101110010111000010001001011011001100001101011101001011111010000101000100000011001011001; 
out3301 = 128'b01110001100011111000100111000011000001010001010101110111010000010000000101010111111001010111001011111001010100001001001111100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3301[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3301, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001101001111110101000001010110100001101010011111011000101010000001101111111010110010000011010001100011001111000100100000111; 
out3302 = 128'b00111110000111011000000001100110010011101010110010101110010011110110010000111110100111101001100011111110100010001100100101011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3302[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3302, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000101000101010101011100110110000100101100101000001101001101110100001001011110111011001001000100011001100011100100111000000111; 
out3303 = 128'b00110111010000001010101000001101011100100111000000100101010010010111110011011100101111010010000010110000110011000101111011000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3303[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3303, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010100101101000011010101110010000101101000010111100010100111101111001000100010000111011011010100011011011111110000100011000; 
out3304 = 128'b11010001100101101010110100011110001101111100101110101100010011100000010111111010110001111101011011100111001100011011001101000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3304[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3304, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101001011101101110101010100100000111110101000000111110101101011101101001111000000110010101010001001010110011101001000011111; 
out3305 = 128'b10100011010000110000111101101010110100010011110110010010101011110011010010010011101000100111001011100100011010101010000011000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3305[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3305, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000100100111010101001001100111011101011101001001111110101010101011110111000010001100010001010001111001111001011101110111101; 
out3306 = 128'b10110110001101110100101010000010100001100111101110011100110011001011110100101110011100101100011101100111000000111100100001100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3306[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3306, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101110110011100101001110001010111001011001101110110100100111101100111110001111010110111100011111010011000010000101111101100; 
out3307 = 128'b10010110011101101010111000110001101100110011011001011100010001110011010000011000000101000000110110111110101000000110110110111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3307[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3307, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000011111100010110011001011011001101001010011100001101101100101011010111101101011101000001001011011110110000000111000100001; 
out3308 = 128'b10000111000111100111110101100011110111101110101111101100001000111011111110111110001101000001001101111100111111001101000110010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3308[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3308, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111010010011001001110000010111011001000111111111100011011000010000110001010101110110000000111101100011001000011101111000100; 
out3309 = 128'b00101010010000101010001001110001101011011010100111101101100100110100001110001010010000001110111010110100011101111011110011110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3309[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3309, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011100010111101111010001101100111110000010011101011110101011101110100110100111101000011100100111101001000011110110001011100; 
out3310 = 128'b10101010000001000011110110111110110111011000110111111001011010011011111100111100011011001011101010011000011101110101110110111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3310[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3310, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100101011000000001010110001000101110011000001100100001110101011101110111011110101001100001110100000110111000010111100011110; 
out3311 = 128'b11101110110001001111101100111000100010110111111100111001101110001011011110010000101100001000001111111011111111101111110110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3311[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3311, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101011100101111110100100111000110001100010010010001001011011111010101110110111000010010111110001100000111011100100110100110; 
out3312 = 128'b11011010011110100011001000111111100101011100110011010011000110000101100011100111101110001000101000111010101001001110111111000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3312[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3312, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011001101001100100000110010010100001000101011010000011110000000101010111010100000101000110011111110010100100001110100000000; 
out3313 = 128'b10010011011000100110111110011011100101001110110010000101111110111110110110100111100010110110001111100101111011100000101110011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3313[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3313, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010000100110000000001110111011110010000100011100001100001011111101010001010101010001100110100011000111011010001110111101110; 
out3314 = 128'b10010011100010111011110101011011110110001100110001110110011111001101001101011010001111100010100001101110110001111110101111010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3314[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3314, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000101000101011011111110010011110001101110110011011010011011100111000000000011110011011011001110110101110010000011000000100; 
out3315 = 128'b10100001011101110100001100101101010010000000101011010111010100110011101011001100110000110000001010011110000000100011001100110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3315[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3315, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001101111000001000011001000100101000101101000100111110000000110100010001100001100001011010101010001001011100000101110100110110; 
out3316 = 128'b10111001110011011001111100001111110011101100001100111000000100010110111101100000111001010111010101011100000111011010000100110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3316[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3316, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110000111000110011010101000111001101101001011111100111011110110000000100101100001001011010010101100010001001111101011011111100; 
out3317 = 128'b00111001101011000010100001111000010110100101011000100111001100101100110000001101111011111100000100001111110011101001001011100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3317[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3317, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011000001000010100111001000100001010111100101101101100000010000111110011010001011110100111110011100111001011101010010010111; 
out3318 = 128'b11000111011000010011100101000001110101010100111100101010100100101100011001011011100011101111100011011001011100001111111001111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3318[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3318, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101111000100100111101100001111110011110110010000100011100000011111100100100101010100000110100011001011110010011100011111011; 
out3319 = 128'b01000000000011100011011100000010100100000110111011101111000000110011100110000100100010110101000001101001001000101010110000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3319[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3319, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001001100011110011000010111011010111001101110110010001000010011001101100111110111110010100010111100100111100010110010011100; 
out3320 = 128'b11110101001110000010101110100110101101110010001001010000111010100001010010101100111101110100111000101011011000100100010100111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3320[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3320, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100110101011011101011010000010101110000110011100110100101100011011111111101011110010101100100110000011001100001011110011000; 
out3321 = 128'b11001011011110010011111111010111101001101000101110101001111101110111100000100011111000000111010010010110101010100001100110100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3321[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3321, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011111111000011101111011100110111011011011010001101101100101001011100001110110001100011000001001011010001101110111110111000101; 
out3322 = 128'b00111101001010001101010001100001111111101100111101001001100000101001000100001010010101011011000101011011101100010000000010111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3322[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3322, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101000001110110010011001111111100011011111000011010111010000001010010000111001110011010101011010000100111011010010111000100; 
out3323 = 128'b00011011100001110001011000000111111100100010110111110010011111010010001100100000011000011111101010111000100000011101100101011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3323[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3323, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110011100001011101100011100110011011011011000001111100010000101000011111001110111000110110000100010001100111001101001111000; 
out3324 = 128'b00001100111010111100100111001010010101100110010110011100000011101010100101110011100111101010101010001100011101011101001011000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3324[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3324, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000010100101001111011001011010111100101011000100110000011000011000011101101110010010111100111110101000101101000011000101000101; 
out3325 = 128'b10110011000001010011100010010110100111111010111101010110011000011100001011011010100110010100001000010010101101010101111111101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3325[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3325, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011111000001000100010101000010100111111011001110001000110101000100100100100110110000010011101101010001100001010010011100011; 
out3326 = 128'b10000110100111000011110010010100101011100011100011101100110001011000001110100110111111010110001000111010110010100100100000100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3326[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3326, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000010110100010001110011110001000111101111000011010111010110001100011101001000010100111011111101000010001100010111011010001; 
out3327 = 128'b10101010000010011100010001110001001010011010111010000011001000001101011100011101100010110111111011000011011010111101101100111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3327[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3327, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111111011101001011001111000101001111001001011110110010100001000010001000101001111011111110001100001101110001001000010001101; 
out3328 = 128'b10101111001001110110110010011100010101110100111011110000010000010011110000000010100010111010001000010100011011010100011111101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3328[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3328, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010000010011000111000000111010000011000100111111110000000001111001001001100001000011111100011010010100001110110101011011101; 
out3329 = 128'b01111110110011111011110011000001101110011101010011111011001001011000001111110001000011111011010000100001101011000100011001000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3329[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3329, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010001000111110100101011110001010111101011111111001110101110101110110001001101101111011000001100010010000010111110010011111111; 
out3330 = 128'b01000111111101000111101000100111010110001100010101010011111101110100100100101111101101110101011000001100000010010101010010011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3330[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3330, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011100101111010010100110001011111011111000000101001111000101100011010101001011010000111010100101011010111001110101011010000; 
out3331 = 128'b11101001010010101101111001010001111111110101010110101110101001111000011110000111011001000100001000001101011111001001101110000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3331[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3331, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101010100001011010111011101110001100110000010110100001000110000110110001000111100111010001001100000101111001100111101010000; 
out3332 = 128'b11101100000101100001001111111011000010000011101010011110001000000001000001110001110010011111001000100101000100100110101000111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3332[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3332, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000001110010000101001001100001111101011011001001001000001110000110010101010101110011101111111100101000000111010110100010001; 
out3333 = 128'b01001010011010101000000000111001111101010001111001001100110110011100101010011111101100000111011000101011010101100000010010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3333[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3333, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100001001110101010100101010010101011111010010001100111101110101101111001010101111111110101110000110100101010010101100001111; 
out3334 = 128'b10010011011001011000010000100010001010101000010011111100011000101010000010100110011000000100101010110101111010010100000100011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3334[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3334, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001100011101000111001110000010100110011110001101001011011000011100010101001001011010010110110100111111110111000011111110010; 
out3335 = 128'b01101000100001110111010100111101110000000100010011101010100011100101000010110000000101011101000000011111011001100010000010011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3335[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3335, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111001100111110011110101110101010101101111111110000000110111111110011001011101110101101100111101000000110001001001010011101; 
out3336 = 128'b11111011001110001011011100101101111110011000111111111011111111001011010011000010011000101111100100111100110010000110111101100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3336[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3336, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010101101101001110100010010100111111001111000100100000000010110000011100101001111011000010001000011011011001001010100011000; 
out3337 = 128'b01110011111011000111010000111100000101101010111001010111111111000100010010000001100111101001011010101100010111000110011011011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3337[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3337, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010011101100100101110101011011010001110100110101001111011110010111001001100100000111000100101000010001111000101000101000110; 
out3338 = 128'b10011101101100001001110000001011011001110110111101001011000001100000001110001111101111000001110101010011001100100100001000000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3338[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3338, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000010011010000100000111100111101010110100000011101000010111010110100101010111001000111111001111000001111110101100001011000; 
out3339 = 128'b01011100110000001010100011101101000101101010000000101101101101011010011111000111011101111100010011100001000010011011001100101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3339[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3339, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100011000100100010000101000001111100110001001010110001100110111010110010110100010101001000100101000000101100101100000000001010; 
out3340 = 128'b01101000000011011010000101000100111001110111000000010011000010000010100001111111011110011011000101011000100110111010101001100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3340[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3340, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111101000010110101101111111000001001101101101011001110110011011000100001011001010001101011101001111010011100001111110101100; 
out3341 = 128'b00000111011001111000011000100001111101000100011011110101101100001010101101011100011100110111001101011011100111010011011101010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3341[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3341, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011010111001111001000001001010010011101000010101101101110011111101001001110011111111001010100001101100011000101001011000001; 
out3342 = 128'b10000000001001010101011011111100110011100110101000111101110100010010010111001011001000101110100110111000001000110010010010011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3342[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3342, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111000110010111101111101101111100011110101011011011011101101110100010010111011100111010101110000001000010010101000010100110; 
out3343 = 128'b11000000001110010011111110000110010111001100111001101010010110011010001001100010110110010010110000000001010010100100111000110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3343[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3343, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100111110001110111011100110100010000101010100101100001111111000011110111001100101010010000011111110001000100001101100101000; 
out3344 = 128'b01110000001101110110100010000010001001110110110101100000100010111100101111000001100100011001000100001010001101110100001001111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3344[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3344, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001111000010101110010011000100010001111100100011011101111100001000011101101001000001101001100000000101111011111101111111110; 
out3345 = 128'b00110011111000111001001110010100001111000110111000000110110101011001000001110000010010000101101011101000000011100010110011001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3345[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3345, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110101111010111100111101010010000011101001111010001010010000001110100110101001111101100110010110101111001101011010001010111; 
out3346 = 128'b10100110110000110100110010101011001101110011110000001001111011011111100111001111000010110100011000110110001100101001011000111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3346[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3346, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111111001011000111001001100111000100010000110001101011011011010111100111001000010011110011101010010000001010100110101011101; 
out3347 = 128'b11110001010001011001101111010011101010011010110000010111001100100101011000010110101100101001100011010010101101010101111110001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3347[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3347, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010001111000101110100100010110001110000001101010011000001001100111100111111001000010011100000000100101111011001111110010011; 
out3348 = 128'b10001011011011111000010111010001000111100001111010010011001010111101100001111011011011011000000011000000100000111011010111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3348[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3348, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010011011001011010001001101111001110101110100001111100010011100010100001111010011001111010110101011110100001010100001000001; 
out3349 = 128'b11100111101000000100001100001000010101111111111001010101111100010110001001110111000000000101001001100001011100100100010011001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3349[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3349, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000010010011101000011110000101000010011100101000000100100000101110010001101001000100101100101001000100001010010000011001010; 
out3350 = 128'b10111100110010011010011011010011100000111000110011110001000000111001010000000110101101000101010111110101011000001001001110010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3350[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3350, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000101100100001010000111101000011101111111111100101000100001101100110111000111111010001011100101001111011101011101010001110101; 
out3351 = 128'b01101101100100000101101000100100110011010110111010101100101000110000001000001011111111001010000101111100101011010001001001111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3351[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3351, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000001000101011000110010010100101101010110011111110101000001011001001001001000111110010001110001101010101011110110011000011; 
out3352 = 128'b00111111000111011100110111101110011000001111100111110010110101011010000100010100110011110011001001100001111111001101110110010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3352[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3352, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110010110011010011001101010100111010000101001000011111000100101000100100100001110010010011110100001111010010010111010111100; 
out3353 = 128'b00110011010000110010010110110011100100001101001010110001101011101101100001111010010111111100010101110000111111101111110101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3353[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3353, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011110100000000100011011111001111101111110110101010110010111110110101101010111101100110010000110100101000011001100101111100; 
out3354 = 128'b00001000111010000111000010110010100001100111010010011000011001010110000001111010010011001001000100010110001010000011111101001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3354[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3354, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100010011011000011101010110001111000011010000001100011110101111101100100111000110101100000101110101010001010110010000011011; 
out3355 = 128'b01011000000000010101010100100110101111001101100000011010111100111011100010010011111100000101110110011000011100101001110100010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3355[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3355, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000100110100001010001010111000100011100011010110100110110001000011001000111001110111001011111010100001100010000010001010110110; 
out3356 = 128'b01000001101111101011101001010110001010110100101110011111011110110110000100111111101010001001010010001110011011101011110101001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3356[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3356, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010101000101100100111110100110001111010101000011101011010100110011011001011001101000010001111100101010100100010110111110101; 
out3357 = 128'b11001110101011010110101000001011011001011011101010001000101010001000011010111101000100111000011101100110110010100010001011101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3357[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3357, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101100101000111100001011000010001110110001000010010110110001000011011101110101000010110000110111011111111111111101101010011; 
out3358 = 128'b00011001011011001010110011011000001101011110010111110000010100111100100000111101101110100010000010011011010110011010100000101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3358[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3358, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001111110010111011010011110011011011000001100110101101011011111001001001101110111001101111001001110001100101100100011100100; 
out3359 = 128'b11001011110010100001110101101101000100010001101111101010111001001001010100111111111111010001101100001010100001110011111101111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3359[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3359, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100100110110110111001001011000111000011001110010010000000011010011000111101100111101110101110001010011101011110111000011110; 
out3360 = 128'b00100101110010000101000000101110010001011100011111001111111100100101101111101101001001011000101110101100000000000111000110100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3360[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3360, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110010101011100101101001111001000000001010010000010001110011111100110110010000000010010111110111001000110011011101110111101; 
out3361 = 128'b00011000010111111110001100100101101001010010000010111110111100000101010101110000000011111111101101101010011110100001000110110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3361[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3361, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101101010000101100111011001001011000111011011001110011011111101110111000011110111101100100111100000010000110000100000101110; 
out3362 = 128'b01001010110100101000100111001001011100110111000110011111100011101111111101011110101000110101110100010100011001111110111100000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3362[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3362, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111110010101110000000001101100100000100010000001101111110000000010001110001001100000110001111111011110111111001111000001111; 
out3363 = 128'b01111111100100111101001001101001110101110011000111000111011011001011110010111011011100000010111111011110000010001011101011111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3363[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3363, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001010100101100111101010110010011110100110001100001100011011111011001000100101100101100110010101101110001100011110100010011110; 
out3364 = 128'b00010111100000000001111101011101101111000100010001100011101101110000000000111000111001010110011011010000101001101111110110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3364[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3364, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101001100000111111110000011000100011011001011111111100110111111111100011100110110110001100011100001100100110100101011100011; 
out3365 = 128'b10011010000101110010101011011011111010001001010100011001010001011001010010011001100111000010000000111011001000101111010100101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3365[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3365, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010010011010110101011101000111111010010111110101000100110001001011000011101100111111001110001010110110101111110000011000110; 
out3366 = 128'b11111010001011100010100000011010001111011000011101010001010101001010100010101111111011011001000101001011110110110010010011101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3366[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3366, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000101101001111101111111011011110000101001110001110110101010001101010010010010001000001000010110000110011110110011011100000; 
out3367 = 128'b00111101000100011110001110110111000001111100011010011110101101000000101011100000010000011100100111100010101110000100000101111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3367[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3367, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101000010111011011011100111110110010111111010110001001011110111101000100010001111110110110110110000111110001101111010000100; 
out3368 = 128'b10000001011010110111111111100001110010111110001101111101011101101110011000000001101000101111011010100110111110011111110111100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3368[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3368, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110010111101000000111010100110111100000000100011000101111001000110001110000101001101110111011001010110111100001011001000111; 
out3369 = 128'b01111111000001100010100100111101000001110000011001101001110111101010101101101111110111011000100000001111001000001100101101110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3369[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3369, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101111000101011101010010011111000010100111011101010111001100011000011111010100001100001001100011000001000101101011110011110; 
out3370 = 128'b00111111000110101100000001000011110000000100000001010100000110001111000110101110100001101001111100000011010111011110010100110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3370[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3370, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001010000011010110011100001011011010110101101010101110011011111110001111111001011000010001100111001000001111101101110111111; 
out3371 = 128'b00111111110010111010000001011111011110111100110000100100100001001101011100110101010001111101100101010000110011110110000100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3371[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3371, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100011000110011100101011010001111101001100011111000110001100011000011100111101111111000101110101000101010110000001101111101; 
out3372 = 128'b11001110100001111100011010000011100010000101101011010011011001111010001111100011101001110111010110110010110101000111011110001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3372[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3372, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110000010110011110010010100111000111011100001100101010110011110110100101011111110100110100101001000101010001110110101000000000; 
out3373 = 128'b00110101111010110001001010011111011111110110011110100111001101101101001101110000001010010101011110010110100010111001110010110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3373[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3373, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100011100010101100001100110111101111110111010101011001011100111111110111110100100010001001100011001011101100011110000101101; 
out3374 = 128'b01011011010100000011011110111010100101000001000100111001011011001011011110110000100111111100111010000011001101101010000101100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3374[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3374, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110111100110011001101010101000100111100010010001110001010101100001010000101100000101010100001111010010100001100110000111110; 
out3375 = 128'b10011101111001101111111000001101101011101100100101001110001001001000111011011011110010101000011011011000001011110001011100010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3375[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3375, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110000110000011101010001010010001100001001100000000111011100100010001001101000000100110001001001010100011100001010101000101; 
out3376 = 128'b11110011001101011011011011111111001111101101100011011000100101000101111001100001011110001110111101010001000000110011110001100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3376[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3376, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111110100110101101000100010101100000000111011100101111101010110011001110010010011000000011110010001100110110111100110011110; 
out3377 = 128'b10001010100110100000001001111010001100000100101111001101111110100010011011101111111110000010111101001010101010011000110111101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3377[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3377, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011000111111110100110011111001111011011010001000011100111110011010100000010110111111000100110001011100101010010010011001111; 
out3378 = 128'b10000100101111010110001001111000110101011110010110001100100010101111001011101101101111011100011001111001010100001011001011001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3378[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3378, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100001111011100000000100011110011110110010110111110101111101100000001011011011111011010110010001100000011110110100100000110; 
out3379 = 128'b10001000110101110001001011100101000111111010000100110100100011000001000010110010111100100111000010011000101110111000000000111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3379[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3379, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110101001111001101010110101101011100110001111100001111010111110011011000011101001000001001101110110011000100110010111111010; 
out3380 = 128'b10110001000101111111000100100101011010010111111110101011000011001110100101001110111100111101111110000011010101110010110010110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3380[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3380, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111101011000100010110111000101001001100010010100000111011110011001110101110000111001000001100101101010011000000010111011001; 
out3381 = 128'b10011011010101011101010110110011101111010010010011011010000001000100011111011100011101100111010011101010010000101011111110110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3381[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3381, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001000111111000110000011001110100011110101011100000010100101101101010110010010111110000011010011101010010100000011001011111111; 
out3382 = 128'b00111011111000010010000111100101110010110100111101011100000000011101011001011101000110100000101101101001101001011100101000111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3382[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3382, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000100010001010111101010000111101100110101010011110000100110001100101000110101000001010101011011010010100111111010100010100; 
out3383 = 128'b01100000011101111010101010110101011101111101100001111011010011101000101010011000110001000101111100010001001001010110110111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3383[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3383, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011101011110001111000110100110111100001001101110100110010110011101010111101110101011110110101110010000101111111010001011110; 
out3384 = 128'b10101111110010101100100001010100011001001101011100101110000100101010011000100011100100111001001111001100011110111111110100110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3384[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3384, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100010000100010101011110010101100011110010111010011010111100010000011010000100001010111101000110101011011111110100000000000; 
out3385 = 128'b00001010110100011110001011101101011011011010100001100001101000111111001100001011111000010101000010100110110111001100111011011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3385[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3385, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011111100001110001101101111111010111001111111010010001001111101110100111111001110100011100111101010101010000000100111011111; 
out3386 = 128'b01000010001000100010111000010101101001111001001100011000110110100111111011001000011110001111100100110110001000000011001100100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3386[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3386, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101101101111000001110100011100101000010100101111100000001100101011001100011010010001110000001111010010101010101011011111111100; 
out3387 = 128'b00111001111011000100101110100011001011101100011010010000101110000010010111001000010010100000001110101010101001100000010100111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3387[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3387, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001010010011001101001110001000010001101000111110101011000101001011011100001111001011011100010111011100111000010111100100110; 
out3388 = 128'b10110111010111100101101110110100011111010001100111110110111100100110111111000111001101011101010111000011100001100110011110110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3388[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3388, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111101011101111000011101110100100101100011001100010110010001101101110110101110101110100110100101100100000001000000110010101; 
out3389 = 128'b00001011100010011000100110111111010010001011000010100110010001010000110110101000101001010011111111110111101101011101111011000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3389[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3389, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110110011101000010100100111000101000111001000110110110011011111000010001001010011000000100111101101110101000100000001111011; 
out3390 = 128'b01111010001110010011011001010101011000101001111111110010000001100010001010101110100001111011001101011000111101111100101100111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3390[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3390, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001111100000111001100101000101110011011011000110110011001111001001100010110110011111100101101110000000111111001010101100100; 
out3391 = 128'b00011000001100100001001110000010110010110001101110100111010000111100000111101110101011110101011100011011100001010000001000101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3391[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3391, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010100000101111011010101101111100011110110010101001001001101011000010101010010000011011101101110001001001101101010010100001; 
out3392 = 128'b01001100001100110011110001000011101100101010111000111011111010001100001110111101001101110111101011111111101111011100001100000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3392[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3392, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101000110100000000000011111100100011111110011001110000010101001011111010011100010011001110011000110011011100000001011000111; 
out3393 = 128'b00100011000110011111010101001100111011101101100100000010001000010100010001001001100001100111111100101110110000000101100000001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3393[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3393, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100010000010110010001101100010010010011111000101111011000101100010001000001011101001111110101011001101000011100101001011101; 
out3394 = 128'b11110010111000011101011101001010111011111110010011110011110010011001100001100000101011110101001010110101011111011000001011100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3394[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3394, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011111010100110100110001011001011000111011110001110001111010000010101011100000011000100001101110100010010010011011110000110; 
out3395 = 128'b11110000100100010111100011111010001111010100001000101110011101000011101000100000110000100101101001111111000011101000110001010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3395[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3395, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110001100111011001011111110101001001111110111001101110001111110011101000000101101110001011000010010101111000010001000011001; 
out3396 = 128'b01011000111000011010110100010001001101011110000000000010111100001110101101000100110110001001010000100111100101110110111000010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3396[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3396, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010101010110011000011001110101111111101000100011111111101001100101111110011010101011101101101010010000011000101101100111011; 
out3397 = 128'b11101101011011110010010001100100001101101010001001001110010001000111111111101001001101001111001011010011001110011101010100110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3397[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3397, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011001110100011100101100110010110110101100011101110101001110001011111100010011010011000010101101110110100001101111001011001; 
out3398 = 128'b00001011110110111000111011001100010111000000100010100001010111101110011000011011101010110110011011011001000000011110010111111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3398[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3398, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110000010111011111110100100100101001100100100011010010001100100001111001010111101011000001101110000001110111111010100101011; 
out3399 = 128'b11111101001000010111001001000000100110111001000111111010001101100100101111011011010110011001111011110001000011001010100101011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3399[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3399, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110100100000001001000000100010111011110100100000111001001110101110110011011000110001000111111101110110101111000011011101011; 
out3400 = 128'b10110000100000011001100010110111011111111001110110001100111000001100000011101111001010001001001010011010101101110010111011001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3400[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3400, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010110010000011111110011010001001111011011111010110000100011010011000110111001000011000101111100100001010110011110111111000; 
out3401 = 128'b01101100110011010001100011010111010110111010000111111000101000111001100111111110011010100000001000101010001100011010010000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3401[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3401, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010111001001101101011010111010001101111100101000000111001000110010100000101001100011100101001100110101110010001101001000100; 
out3402 = 128'b00011010011010000110001111100001111011100100010110001110011111001010101101000000110100110010011110000001101001000101101001111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3402[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3402, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011110100001111111001010001101010001100010001011110011101110101100100011001100100111100000111011001010101100101110111110011; 
out3403 = 128'b01011001110010100101000000000111011000100010000011001001111001000111000001000010000011000110011111111100110100111011110010001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3403[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3403, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011101010101110000011100000010001011000101010010011001001110101110000010110001111011111110001010011111101011000110011001111; 
out3404 = 128'b00011010101000111100101100010010010000000001010100001101110011010010010101000001011011101001111110100111101010111011101100000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3404[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3404, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011000101001111011011100010011110001011011101010101101110111100010101111101010011001010010111001101110010100000111011100001; 
out3405 = 128'b00111101000100111101001000000000011001001011010000010000101100101111001111001101011101111010001101110000000000111001011010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3405[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3405, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111001111011000011001000100101101011001011110011100100111101101010000000010000001001100101011100100001100101101010100100001; 
out3406 = 128'b11001010011011001000100100111000111000111011110110010011100010011001011110101011111110001100101011111100000101000111011011010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3406[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3406, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011011011010011101111010100011110000100111100111011100101000000001011110101101111110001101000110011000010100110001011011011; 
out3407 = 128'b11000000001010010111010101011011011011000111110101010100100101000100010011000100001001110101001011110011111110110100110010010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3407[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3407, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000000000101101111001010110111001010100001111101101001011101001001101010110100000000000000110011110011101100000100110001011; 
out3408 = 128'b11111101010001100001101010001000100001010000100000101001001001101010111011101001111100100100110000101100110100111010110011001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3408[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3408, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010110110010010010100101100111000010011011001110001001010100101110010111110011000000010101100101001100101000011000100111011010; 
out3409 = 128'b11000110001111001110111111000111100001111011110101000010101100100111111000001111110010111110111111111001000101001011010100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3409[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3409, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101100101111001011100110100101110010101010101011100111010011001010100110101001001000111111110110100111101001100111110001000; 
out3410 = 128'b10001100010001010100101000111100011001101111010101000010001000011001111100111010110110010100010011000100111111100001000000101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3410[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3410, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011000111010010010110111111010101010111011001011001100110100011101101111111110100011110111011110000011011100000001010001111; 
out3411 = 128'b10001110000000011101001111110001001111000100011000111111111101101110100001101110101101001000000111110111101101111101110101010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3411[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3411, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000001110001101110100111111110001111101001110010001110011000011110101111110010110010000001101010100000110111010110001011110; 
out3412 = 128'b01101010010001000110000000011000111011111111001101000001001001100010001010111110110111111111101100001110011111011001110111001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3412[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3412, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000100100100011111110101101000000000011101011001100011000110110110110110000110000001001000001010001000001010011101000011000; 
out3413 = 128'b10001110101100110010101101100010110110111101101000011100011010101000110011111011100001010010110100100111000110011100011010101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3413[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3413, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100100101000011000100111001001101101001000111101011011111001100000010101000010001110011101011100000010101101110001101111100; 
out3414 = 128'b00001100110101001011101111001101010000000000101101010111100000111101000011111110110110110111111001001100011001110000101000111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3414[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3414, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000111000001111000101010000110000111111000001010101001000111001100111101010010011100110101000101000100010001010110011100010; 
out3415 = 128'b11011000001010000100100000100010011000000010110111111000101101000100010111100101000010010011110110000000000101001101100100110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3415[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3415, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011110101111100010110000011000000100100001101100010010111011000110000101011111010011000011100101111111011001101010110111010; 
out3416 = 128'b10010001011111000000111001000010000111001011101110001000111010010001010100101011010101111000001000111001110011000010011100110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3416[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3416, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101110110100110111101100010001111011100001000111101011010010001111101000001001001011000000111010010110000000111010000001011; 
out3417 = 128'b10000110011011001010010010001010111010100010111001010010100111001101100101011111001101100101010110101100101111010001011111011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3417[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3417, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111011000011001101110011100100110110111101101110001100010101111001100001001000100111010110101001110100000111111000001100011; 
out3418 = 128'b10011101010011100001100000000110010100101100101001101101001110110111011101100110101100100110000000100011000110110101110101011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3418[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3418, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010000011000001000101011101100000100001111110000001001110010001001110001111110111110111110101011101011000000001001110111110; 
out3419 = 128'b10100001000000000111111100001001000001110110010011000110101001000110011110001101101010101100100111011011010101000011110010111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3419[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3419, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010001110101011111010110111010101110000100100000010000011110111000101101100000010001100110011111001100011001111010011100111111; 
out3420 = 128'b10010001011000000111100101010001111001010011001000000000001100011111110110100011010001101001100001001010101001100010110011110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3420[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3420, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111100111110100010100110001010110001101100000001001110011011111111101111110111100100010000100001010010010101000111100101100; 
out3421 = 128'b01100101011000010001110110110110011111010000001101001000010110100000010010000011100010110110001100100010110001101000100111111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3421[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3421, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001100000100011010111010110101010101110111100001000110000101111100110101010100011101011001001010011011011001000010001101110; 
out3422 = 128'b01110110100011001100110011001111010101110101111110110100101111000101000010001011101110010010111100111001011101001011101011110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3422[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3422, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111101110011110100001010101000001011111111000110111111101111010011101010111010110010111110001011100000011101100111000011011; 
out3423 = 128'b01111000000001101100110011000101100001000110110111110000101000001000111001000101100000010001111100111000110100101100001101110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3423[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3423, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010010110011100010100100100110110010101011110001011100001000000101101111010000000000001110101001111111000010010100111001110; 
out3424 = 128'b11001111100100010011000000010110011000011010111100110011101101100000110011100011001000100100001100001110011000110110010111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3424[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3424, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010001000011100111111011010111000000000100000111000001111101111010011001001001010111000101111111100000110110011011001101110; 
out3425 = 128'b00000110001001101000010000110110111001011000111001010100010101111110010111000101101001101011011100101000011110101011101000000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3425[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3425, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110110011111000111101100100100000101111001001001101110111100110001110011011001111111000101011011100011110000110000110001000; 
out3426 = 128'b01110001010000010000100111110010100100001111101000111000010001011100111110111111100010001100000111010111011011100111101011111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3426[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3426, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111100001010010000100100010101011110001111000100101111111110010011111001010010110000101101100000000000110101100101000111011; 
out3427 = 128'b00101010111000100011010101011101010101111110110111111111110011000101110111000111100010011010111110001100101110101000101000101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3427[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3427, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001011010110011010011111110111000111111110010010000010111001110010110010110101111011110101011000011000101010100101110100100; 
out3428 = 128'b00000000010010111110010101110100100101100101000011111010101000000101000110011010010111010000101110011000110111101101100000101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3428[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3428, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111110001010001000110000000110101111010010010100111110101010100000100110101101111010011011011101000100000100110111100100111; 
out3429 = 128'b00100000001110100110111011011011000110000010010110100101100110000101000011110010111111111111001010011011011000100110111111111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3429[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3429, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001110100100111100111111111111110110110001011101100100011111010111001100011110011001110110101111111011011111001110100011110; 
out3430 = 128'b01011101011011001010101011001010001101011101001010010001001111111000011110101000101000001011010110110100100000000001010000111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3430[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3430, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110000111100101000000000001010101001001010110000000001111010001110001101011001100011101110111110001010010100101100110000111; 
out3431 = 128'b10110010001111100000011001001101110011001100111111101010000100100100001111110001010100111100011101010011110011111111010101000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3431[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3431, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101011010011011110100010001011001101111011101100010010100110011110000000010100011100111000111101011101001011001001101010010; 
out3432 = 128'b10101010000101011110100101001100011111011011000100100000001101110101110011001011100100011101000000111010001011010011011010101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3432[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3432, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011101011011101010011000100000011111110000000011110001100111100100010100000110101011111001001010100011011111100100100100001; 
out3433 = 128'b10110100101011000010000001011000011101110010010001110100001111101111111000110111111101110110010011100010011111001101101100010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3433[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3433, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101111111111101010010111101001001000000111111101100110011000010001001111010100010100111001100001100100110101000100101111000; 
out3434 = 128'b10001100011111011101100110100010101100011010010011000010111111100010011110001100011000101010101010001111001101011100101001000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3434[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3434, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100011010001111110110110101110011001010101111100011100110011010001000011101001011100010010110011010110010000101101010000001; 
out3435 = 128'b11110000001110110100100110100110011100011010001101011000000001010000111110101100011010101000111000010100100111110111010111010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3435[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3435, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101100000011010000001000000010011110001011011100101111010110110010011111110110100000100011111011000011100010001111101110101; 
out3436 = 128'b00101001000110100001110011111100001110101110011010000110110011110100111111100011001100011110001010000001001100100111011001001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3436[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3436, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010000100001001011111101011111010111101110010111101101111001111111101000001111110110111011111010111101000011101111110010101; 
out3437 = 128'b11001010010001010001010011001011110100010011010101000010101110111001110001100000011001101111101000101000111001001011011111100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3437[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3437, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100001111101000000010101111100011011100111101111010111111101010111100111010111010001011001000011100100011001111111010101111; 
out3438 = 128'b01111010010000100111100011001110001110001011010110000110111000010110011010000001011110111001111011111011100110100111101001111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3438[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3438, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110011011001111001010011110001111010110110101010101000011101110000100010001000011101010101111000101100100101000110111000010; 
out3439 = 128'b00111101010111111011101010011101101011101010101111101001010111010100100010001010000101111101010111110110111101000111101000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3439[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3439, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100100110010000111100100111110100010001101110100110101000001001010011001010000100100101001011100110011011101000101101000110; 
out3440 = 128'b00010110101000011101010010110001110100101001001100011110000001001011110110110101101110000101010101011101110011010111101001001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3440[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3440, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100100010001100011101001000110111000001010100000001111101000000100011110000001101011101010110011110000001001111110010101110; 
out3441 = 128'b11100010100011111001101010001011111101010011110000001011111011101101000111100000011111010100101010101111100101011110010101011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3441[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3441, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011100000111100100000110000101001011000000111101001111100110011001100010111101001010001101001000110101011100010000111101111; 
out3442 = 128'b11111110001111100101111100011001010111100100110000001110000000100101001010001100101010101001011101010111101011011110011011111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3442[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3442, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000000110000111011000001011100111000010100101000001101000110100101011111100100001101111000110000001111010011111100100001111; 
out3443 = 128'b00100000001101010011010110011110110011111111010101101111101010101010001110100000000010010100111001010110011110011000010001100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3443[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3443, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100011100011100100010000101001110011100110011110010010110111011100101001111101111011100100110010110001000001111100101111111; 
out3444 = 128'b00111011010011000010001110001100111100010100000011011010101010010100011110110011001001011010011110100010001000100111101001000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3444[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3444, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111001001101011100100001011110001100101000010111111010100011011010100000100010111110111010111110111101101111111000011110011101; 
out3445 = 128'b10001100010101011100100111010111111001101111000100110100011001110000100110011101101000000110111000010010111110110000010010011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3445[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3445, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110001100111100011011110101011010111010000101110111001100111100011101100011011111011010010110101101100100111101100001000111; 
out3446 = 128'b10111100011111011100111100110001010101010111111100011011011100110101001101001101011111011110101001101011010010000100111000010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3446[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3446, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101101000100010001100110011101001110101100001000010001101001111001001011010010011110101011010101111111001110110011100100110; 
out3447 = 128'b00010000101101010011000111100010001100111010000011010100110001100110100111100001111011011010101111000000010011111010000010110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3447[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3447, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000011001001011110001001010100000110111110101001011111100110100011011101111101010010111101010010011011111001001100001100010; 
out3448 = 128'b11111100011001101011000101011100111000100101111010010000001100110111100111010101111100111001000110011010001000000100000111100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3448[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3448, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100001101011111101010100000110000110010111111000101011000101110000111101011000011110010000001011010001101101011110110010100; 
out3449 = 128'b10100111100011100011111000000100110010011000000010011100011001111010010101101110000001100100111100100110001110010101111110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3449[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3449, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110011100010100010001000101011100100010101110110010100110010111100100100001001101100010011000101100110101101010110001011000; 
out3450 = 128'b01010001011011011110111100111111100001001011101011111001100011100111000011110001111000010000010011010110010110100100111011000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3450[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3450, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000000010011101001110101000101100001101000010001101100001101111101010001101000011001110111110010010101101100010000000011010111; 
out3451 = 128'b00000011011010100011000110000110000000011111101010101000100100101100010001101001111001011100010110010111010101100000101001011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3451[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3451, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001011000000001101001111111001100101101100001111110111011000101001001000011000111110010010000000111001011010100000110000000; 
out3452 = 128'b11100110110000010101001100001000101011001110100001000001100101011001011010010110000011000001001110101010101010001101001000100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3452[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3452, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010000110101110000100011000111100110000110110000001011001101111111101101111101101101110101110000110110000111110011111111111; 
out3453 = 128'b11001111100100111001010001111010111010011101010101100010101101101100000111111011111100111101111110000000011011101100100101110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3453[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3453, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110101011100101000011001010100110100110100010001111100100010110111111110010000111010000011101111100001111001110010110010101; 
out3454 = 128'b00100001100101011100111010011000011110011110110100100111000110110001111000000110001001011001010011010000000001111001011011001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3454[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3454, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101001010101110000001000001101100100000110011001100011100110010001111000111000000000010100110010101100110110001010111011000; 
out3455 = 128'b00101010010001000101111110011110100001010010011010100110010010110100110011011101000110001011101101101111010010011100011001001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3455[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3455, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100110101001110100111110110100001001010100010000111011111110110010000100110010100000001001111101001101010110110100101110001; 
out3456 = 128'b01001101100101001000100001100010110101111110110111101111010011001111000011110111010011111011110000000000001110010000110001000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3456[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3456, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110010001100111101000000011100101100000101101011000100100100000110110001100000010110100100111011101010010110000101111101111; 
out3457 = 128'b11101111010111011101010100000110011100101100000011111111111001011100010100111100101101010000110111001000000000010111110000110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3457[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3457, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100001110100100110100011110100101001111001001101001101001000011000110101100011110000100100001000011010110000100110011100000; 
out3458 = 128'b01101111111111000001111011110101011100101111101101010010010111111100111010011101011111001100101010000111000011001100001100110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3458[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3458, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111001000110011011001000011011010100101001000101111011101111011100010110000001001110001100110000111001010010000011100000111; 
out3459 = 128'b10101010010011100011010111010101010000101011110101111010001111110000000000011010110001011001111001111011100010010111100101111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3459[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3459, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001010011111000001110110101001111100100101110101100011101001011100110010010000010000111101100100100000100110110110000011011; 
out3460 = 128'b10001111000111111011111111000001011010010000001110000100011010111010000110010001101011101101101001100111111101100111001101011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3460[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3460, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011010001100111110110000101000101100010111101100111011100101010010100000001101111100011110011010100110110011001101000111000; 
out3461 = 128'b10001001001111011111100001110011111100110111001000010100100000011010011001010100011001101101011100011011010100011100100110111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3461[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3461, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110100011001110011010111011101011101011011011110100111001110011111000100101101001111001000000010011110000101100101101101100; 
out3462 = 128'b10001000011111110111111000111101000100101101010100010111111001100100100001010111001011000100010100110010100000010011111101010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3462[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3462, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111010000111111010010101000011110110010100100010001011100001100100000101010010101000000100100100110011111100001101001001000010; 
out3463 = 128'b10010010100001000011010110110101010101011100101000000100000011111111000100111011010010100101011111111001000111100101101111011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3463[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3463, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000000000010110110110010101111000000100111000001000100010011000101100001111101101101100001011011110111000101101000111110000; 
out3464 = 128'b11010101000111011001100111001101000110110001110010110000101110101110101000101011011000011100011011001101010110011001100010011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3464[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3464, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010111101100111010100010101110111001111001000110001010101011010100001001100110100100111100001001111001100110010011011100011; 
out3465 = 128'b01110101011101001001110100000111101101111010011110010100110011101001110101000001101100100010110001111000010010111100011100100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3465[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3465, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000111110011011101100100110001100010100111100110111011001111111111100000011101000000001011110000111110110110110011100100011; 
out3466 = 128'b01001101110011101010000100110011110100001010000010100101111011101110110001001111110001110001100110001010101000001001101001011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3466[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3466, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001111110100111110010011100011000111110011010111100000010101111010100010110010001000001011101110001100111101101010111011100; 
out3467 = 128'b10001111100001100011100100000000010110011011001010000001110100000111001100100011011011001101100011101011111111100101100001000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3467[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3467, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001001001001101000011100000101111101011101110100010100001011010100011101010011110100100000111011110000010110101000110011000; 
out3468 = 128'b00011101001111000000010100111001010100111101100010000111101110000011011100101000100000011000101000111010010110110010101011000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3468[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3468, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001010010011110101100111011011100010001000110011100111100000101010001101001100000001110000111111101011100101001001010001000; 
out3469 = 128'b10000001010100101110100001000101100010111000100101100101010111111001110100010011100111010001110001101101110110110110110100101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3469[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3469, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001000001000110010101111111000011011111011010110011001010011000111000100110101101110011001011011110111000010110001010100010; 
out3470 = 128'b01101111010111011001010100000010100010011111000001101100011111101101011000101011000111100001000110110101101010100010111100000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3470[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3470, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100000010011010100011011110011001110001100010101100110100101110011010111000111001110001100111001001011011001111100110100000; 
out3471 = 128'b11010010110101010011001011100001111111011111101001010101101000010011100100100100100000011001000001110101011100000101101010000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3471[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3471, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110001011110001100110100010001101111001011000000101000100101010110110101101111000000010110110001110011111101011101110001101; 
out3472 = 128'b10100011011111110010010110100100110010011010011011000111001001111100110100011001110011011111100101001110100100100111111100011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3472[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3472, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101010110000000111000011000001001100010111101101111101101100000101000011101001011011010101101101101110111011011000010110000; 
out3473 = 128'b01110011110001101001110101101010100111001010010111010101101111000101001001001000011110101110110100110010110110000101101101000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3473[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3473, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100011011100010001000010000100000000100011010100100000110101001001111010111110110001011001010000011010101010001000100100001; 
out3474 = 128'b01001101001011110000000100100001111101100111001001011001100011010011101101110100111110101101110010110100101110001111000110101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3474[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3474, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010011000001000111000101111101101100101011111100110001110010101000010110111010000000101111011101000001101010110101001110101101; 
out3475 = 128'b11010111110010010100000110010110010101011101001101100110111000011011100100010100101110101001001010101010101011001000011001100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3475[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3475, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011110101111001010110111001000010110100010110000101101001111101000110001110111010000001101101111111011001010100100010111010; 
out3476 = 128'b01001100011001011101110110001000111011110000110000100101000100011000011101110011111000100110010000010011000110011101100011010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3476[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3476, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011111010001111100100110111111101101101111111111101100100000001011101011010011101111010000111100001011100000001111111010000; 
out3477 = 128'b10100100100001100100111100111111111111010010010111101100100111010010011111100011010110001101000010010011000001101011111110101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3477[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3477, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001010100111010100110101010111010011011010010011100100010101011001111010000111000111010011011001010010111011110011011010111; 
out3478 = 128'b10110110101010110010001010111000010111001000100010100010101111010111110010100101101101001000001000000000000110101010111101101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3478[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3478, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100010110000100100100010100110010101001001000100111001010001101001001110010000101001101101100000011010011010101110001110100100; 
out3479 = 128'b10101001111101011101010111111010100011000111001000111011110110011111011000010010001001100011001011110110000101011101001100001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3479[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3479, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011011010000110000111100000100010000110000000110101111000010100101011001110100000111000101111001110000000100011001110001111; 
out3480 = 128'b10101111110111110100001110100101011010100101001111110001110000111001001000101110100000110011100110000000111010100111010111010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3480[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3480, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101001111001010101101010001111111001100110111110000000001000001001010011111101101100111111101110100001110111101100011101101; 
out3481 = 128'b01010010101111010011011110110010010010011100001000001000110110010101011110100010011111011111010110011110101001001001111010101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3481[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3481, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111100110110001000100111000001001100111000110000100111110100111000100010111101010001010000010010100100011111001111101011000; 
out3482 = 128'b11101110000001000001010001101000000010100010000011101010110001000100100100001010111100010101010111101011010010010111111110101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3482[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3482, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010011100001111100001001010111111000010001111010000000000110100101011110001001110100010010000111110000111001100100000100100; 
out3483 = 128'b00010111101001001000000010011110101001100000011000101011110110110100001001100101100000110101111000101011011110100010010101001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3483[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3483, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000111100011000100111000111100110101010001001111111010001110100101100110001010011000001110011001010001010100000101010101111000; 
out3484 = 128'b01110000000011111110110001110111100001111011001111010000100111111100011110011110011101110001101001001010101100111000110100101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3484[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3484, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100111110101110101110010000001010110000001100001101011011001010010110000110000001001100111001010000110000010101001100101011; 
out3485 = 128'b00001011101001010001110011110010000110000001111101101001101001001100000110110011111100100101010010011010111001110000111101001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3485[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3485, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100000011111110110101110110100110101010111001101010000111000100010110100110111010110011011111110010000110001110101001100000; 
out3486 = 128'b10010011110001001101011000001010111111000011001101100000000111101001000010000001110101001010100001110111111100110010001001100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3486[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3486, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011111010010101011011001011010001011011001110000101010111010111100111001111110110100100011001010010100111010101100010100111; 
out3487 = 128'b11111100100011011101010101111010111100110101001001000111010110111100100010000100100111001001101010110000110000010010011111111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3487[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3487, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111011001000011010100111111100110111011101011010001100011001001000011110011010111101110001011100011111011010101001110101010; 
out3488 = 128'b01010001111101001101100010111011101001101011001000100100110011000011010010111110011111001000101001000010111000100101010000110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3488[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3488, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001000001011100000111110111010110110101111110011000000110100001111011111101011100010100000011110011101011100111100001100011; 
out3489 = 128'b10000111101110010000000111011010110001000110110110100100101001000000100001111011110110010010010000110101110101001111101100010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3489[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3489, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100100100110011100111010011000110110101001000100010101100011001100010011011111101101111101001101010001111100010101111100011; 
out3490 = 128'b01010001001011001011001011111011101011010001000111101001011100010001110011001100011111110101100010111001000011010011110111110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3490[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3490, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000100000001101110110001010000110000011101010011011101100000110001110000110110110110101010101011000100001011010000001111011; 
out3491 = 128'b11001001110111010101011100000000011101000011000010101110010000111101100000111010000110011000100110011101010011100000101010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3491[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3491, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111100110100010110000001000101010110001010110001001000100010110101000010100101110110001011011000100010110111110010010110101; 
out3492 = 128'b00101100000100011100101111100110010111110100000110111111110111101000100000111111101111011010010101100111011001011001101111111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3492[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3492, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000000100101110111011001000111010110010000000010110111010010101100111010000000100000111101110001010001001000101100010100000; 
out3493 = 128'b01100110110010001110101000111001010011001101000001011010111011110000110111010001111111011011010011100110111101100101110100100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3493[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3493, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111101101111001001001111110110010110001010111011111010101000001010000110101010011011110000000100001001010110010111011011111; 
out3494 = 128'b10111101111101001101011101011111111111100010000111010000110101111010100101000111101011001010110000000011110001111111101001011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3494[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3494, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101110110000111011110011100100001110000110101110101010001001101101001000110010001000011110001000111110001010110010101110100; 
out3495 = 128'b00100111111000011110101101010001101111000001000001010010010111000001011110101010000000111000011001010101010101000001000110100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3495[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3495, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000001110001110001001101011000100100010111010011110011110100000001100101010010101000001101011000110001011010011100110100001; 
out3496 = 128'b01001100111101110111101110100000010111111000101011100010001011101110010100110001001000100010001000111011010010100100001101010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3496[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3496, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100011110000111001101011010101000101011011111101100001001001100000010010011010101101111011100010101010100100111100101001010; 
out3497 = 128'b10110101010100101000010000001010001111111111100111000100111100110010110100001010100100101111010110010001000001001110000101110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3497[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3497, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001111101110000111010010111011110000110000010101110110100011101010111101000110010100101110101011110111111010100111011101101; 
out3498 = 128'b01001111001101101000001001101000001100010001011111100001001100110011100100101101110110111011111011111110000010100101011011100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3498[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3498, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010010100000100011011111100101001000011101110101000111111011011001101011010000101101111011000011011100100111011001111011101001; 
out3499 = 128'b11101000000100111111001100010010000101011100101010100110010001001101011101000111110101110111110100101001010111100101011011011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3499[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3499, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011000111011011101011000011111000011011110000000001010101101000101100110011100110000110110110000100001101101010001101110001; 
out3500 = 128'b11110010010110110001101100100011000110001101110100110111000101011001101010100000101110010001100011001110000110100101110001111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3500[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3500, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000101011111100100101110000010101110101101111111111011111101101100010001110011011001100011000110111010001101110000110010001; 
out3501 = 128'b10010011011101001111010101111001000001110110111100000110010101011111001101000100110100111000100000010001000110101001011001111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3501[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3501, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011110110101101111111001100110001101011000111101111000110101011110011001100010011110101100110100001101001010010111101100100; 
out3502 = 128'b11111010010000100010001111011000000011110011110000011111011101101010100100011101100111101101000100001101011000110101111010101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3502[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3502, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000100000110011000100000000101110111010011100011110001110100000010100010001011100111100010101001110111111110101001111001000; 
out3503 = 128'b01011110110110101000100011101111011000101011111111000101001100100011001010100101010011000000011011001110111101001101000111110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3503[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3503, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101100101011101000000000001100011101110001111001011111010000001000111010001101011010101110001010100101011101010011011011010; 
out3504 = 128'b10100010111101001000110111101011100111000011010101100001101111011000100000100110100011000001101000110000011010100000100100010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3504[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3504, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110011101111111101001011001011011101001001010000011000001001110011011011101000100111000101101101101001001110111001001001111; 
out3505 = 128'b00111010110011110110010000001010101001011000011101000101010101100110001000101011100011010100111011111101001000000010000001011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3505[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3505, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100011101010100101100100111011000010000110100101000111101101010000101110010111111101011101000100110010010001001100101110000; 
out3506 = 128'b00111011001010101000110011011111111011100010001001110110010001010011010010011011001010010001011100110111011110000000101010110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3506[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3506, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110001010110010100000111111001001011100010100110111000100011111000010110010111100111010001011100111110010001011111001010011; 
out3507 = 128'b00000110101001101111101001010101111111111010100001001001101100000110010100000010011010111011110100100101011001010001011001010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3507[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3507, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011001110000100111100101011001010000110010000111010011001001010000101010110000000101110110011001111011100100011001010111000; 
out3508 = 128'b11110101111110000111010000101101010110101110100100010000101101010001000011100110001101001101011010111101111010101111010100101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3508[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3508, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100101000000101000011101000111011111001011011010001100110100110001101001000101110101111101011011010110011111101110011010110; 
out3509 = 128'b01111001111000100000101000010010100011101110010000010100110111100000111001001011101000010111110000111001001111100000111000011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3509[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3509, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110110000101101010001001110111001100001001110101001010010101010010110001000010100000100110001101110110111111010011011010001; 
out3510 = 128'b01100110001110001100010110001011111000110011001111111000110110110000011100111101100010111110010101111101000111111110010011001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3510[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3510, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110001001010010110111100010110011001010000011011010011010001100010110101010101011010000100010100101010101001001101011001011; 
out3511 = 128'b10000000001000001100000111011001100100010010110101000100110011100110110100000111001000110110111101101110101010010001001000101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3511[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3511, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101110101011111111010000111110111011110110001110100100111001111100001011100111110010111101001100011100001110111101010101101; 
out3512 = 128'b11100100100011011000110001101101111100010110011111110001110100000001100010111100101011000001000000110010011100101111000011110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3512[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3512, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110011001100101101001010111001111100111101011011101001101011110110100100011100110000001100100100011001100000110011100110111; 
out3513 = 128'b10011010000100001101110000101011010010101101010011100001111101100110100001011001011100010011110001011111111010111110001101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3513[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3513, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011011100101010100011100011010001001110010010000011011001000110001101110111100100110110010110000000010110010011111101101100; 
out3514 = 128'b01111010100101001001101101111110010110010111101001101101011100100000101101000101111000101100101011111111110011110111111011001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3514[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3514, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011000001000111101011110011000111110111001110001101111001010110111101101001101110010100110010011111010000001010010011001000; 
out3515 = 128'b11011001101010011110010101100111110011110100111111011010110001100001011011110101010101101010000000100000110011101101011101010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3515[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3515, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101100001011111011101100001000010010001100110001010001011110011000001101000101001101000000001100100111100011110000101110101; 
out3516 = 128'b00000101000100000010100101000111010101000111111000001001111110111001110101100001011101100101010010001011101110001100011000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3516[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3516, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110101010000001001010101101001001001111011001001101011001101010100010000010010100011101111000111111111000011110110110000111; 
out3517 = 128'b00010111101011111101100100011111100001011100111100110100011110100101101111000100100110100111001001001100100110111000111001000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3517[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3517, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110001111011101111110100100011011100111100110001010110000100101001110011110100001010111000100111101101001100011111011011000; 
out3518 = 128'b10111111010011100011110001011100010011100110111010110101000010110011101111111111111100111010111001101110100001101010011010010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3518[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3518, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010110110001110110110111011110010111001100110010100100011110001001001101101100000011010100100101001101100000101011110100001; 
out3519 = 128'b00111011001111100010001110111100101010111011011010010010100010011110000101100100001101110001001100010011001101100110001000110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3519[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3519, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010100101000110010100010000101000011110101111100110110000001111011101010101110100101101111010110111001100000101111111000000011; 
out3520 = 128'b10000011011111101100110101110010111000001011111000010011100100000100010101001001000000101000011110110001000011100110101101010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3520[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3520, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010000100111101111100110101111111111110110000000000110010110000010010111011000001010110100000000001011100110010110001100000; 
out3521 = 128'b01011110111010111110011000111111010011110101101000011100011111011011010010101000000110011111110111000111110101110110110001100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3521[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3521, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001011111000000101000001010111111001101011011101101111100100010001011100000000110011111001110001010111000011000001100100010; 
out3522 = 128'b11101101110010111101101001011010000100101001000010011111000001000110001100011010110001111101010110101000100111101110011100001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3522[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3522, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111001111000000011010101011011010000010100101111010001011111110100010110110110110110000100010110011100111100011101011000010; 
out3523 = 128'b01011001011000100110011110011011011000000111111010111010111010011011010001000111011010111001000000101000010101010101100111100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3523[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3523, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110000011010110111100010001101111010010101110000100000000000011000110101101111001000001110010001100110010000110011010010010; 
out3524 = 128'b00101110010111001101101110001010000001010111010010101101011101101100011101010010000100011100011001011010100111111101101100011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3524[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3524, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000100111010001000000010101100101100001100011111001001011111011011011010101110000101000111011101000110001111111001000100100101; 
out3525 = 128'b00010110000010110101011101101011101001010001101111000110110111000100101001111011010000000011000100001101101101001110101101011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3525[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3525, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011101101111001110101110010001010101110001101001011101100001111111010100001101011010011010011101011011000110001111101101111; 
out3526 = 128'b00111011000000011111111000100000100101001011101100011011111100001110010100100100011101010111100101001001010100001111000001101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3526[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3526, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011000110101000110000111011111000010001001101100010100101100000000011011110000000001000011110100011001001010010001100000110; 
out3527 = 128'b10101000011110100110111011001100010111101011011101001010111111001110011101000000111101110010011100011010111010010001000001101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3527[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3527, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000010000100011100110100010010110001100000110001101111011011000101001110100110100101110010001000110011111100110100111111100; 
out3528 = 128'b11101000100101010011000011011000111001110111011001111100110100101010111000101111010101010111001111110000010110010110110101111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3528[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3528, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010100010110100101101000001101101111110000010100000101100001010101100011101010100111011001101110110001001000001100101111011; 
out3529 = 128'b00011011010010101100100010101110010000100011101010010110111011111110001001111100010100110011011101101100101111100101000010001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3529[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3529, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110010100100011110001011011100010011101000101111000010101001010011110111000101011100000000110000010101001001101111111101100; 
out3530 = 128'b01111100110010010001000010110000010000100111100000100100010001001110010111110100001001111011010101110111101001110101000101001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3530[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3530, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111000000010001101100110100100011000010011110111001010000010010110111110010101010101100010110000011100101011111000000001101; 
out3531 = 128'b00011000101011111111110110101100010000000110110000111000110110001000110111111100101001101101111110001011010001010010010111110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3531[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3531, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110000001001010000001001010101000110100110110100010010100000101001011100101111001111111001100010101101010011001111101100011000; 
out3532 = 128'b11010000101010001011000110110101100100000101001110110000110100010111010001010011000000010001110010110100111000100111110101110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3532[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3532, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010101010100001011101100110110011100100111001001011101011001010000000110011010000001110100010101101110011110000111101100000; 
out3533 = 128'b01101001111100000011011001110000111001000000011011000110011110010100010010000001101010000011100000100001111101010100110110010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3533[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3533, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000000011101111111100111010111011100101100111000010000100011110000110110111110111111001001101100111000110000100100010011001; 
out3534 = 128'b11101111100001010100100100111100010000000010000101001101100101001100000010101000010100100101101010110110110101000011110100010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3534[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3534, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000011111001101000110110000110110001011110011100010100110011000000110011101000111110011010111000011101110111110011100000010; 
out3535 = 128'b10100110010010010101000000010110010000110110110110101011011000101010110111011010000000000101110011011011000011110010011010000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3535[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3535, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111100101101001101101100110100100011000101001110111110100100101101011001000111001011111110010011101011101011111010001010111; 
out3536 = 128'b11011110010101010001000110100001100011100110000100001100110000001001000101001100111110111110101111000001110111111110110111011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3536[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3536, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010111001000110111000101000010000101111000001100000101011101001000100000100011001001101000000000100111111111001110100001010; 
out3537 = 128'b10111010010100111010000000001010000011011000010001110111010100101010011101101111110001001000100110100110100111100010111111011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3537[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3537, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011101000010111001010100001001100110111011100010011111011010111101111100100100011000110000110111100101010111100111111001110; 
out3538 = 128'b11001000101100110101011100110001001101110100100011100101000010100001101011011001010100011000110010110010110000000010101011110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3538[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3538, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110000101101101110101000010100100111011011110101000110010001111011100000000010100110010010011000110000110100000011010111100110; 
out3539 = 128'b11011011111010101010100101010011100011001101110001100010100101001111100101011010010110010110011011000011100010000100101101110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3539[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3539, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011010111100000011101100000001101010111000000111011010000100101010010001110001001011011101100111101011001011001001010110100110; 
out3540 = 128'b11100001011000011000100111110101110101010111100110101100111010100100100111000100111100000000110011111010001110000110001100111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3540[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3540, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100010010111111111000010110101110001101110010110110010000011101000111010110001100011011101001110000010001110000101111010110; 
out3541 = 128'b10001110111111001000110101010101010000011111110110010000111000100110001001111101111101110111001011100000111000010001001110000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3541[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3541, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101101000100000011010101000101100101111010011111100000110101110110011110011011111000111011110001110111001011111001101011110110; 
out3542 = 128'b11000111011101011111011101000100000100101010101001010100000010001010100110000001000110111000100101111101100110110111110110110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3542[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3542, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110110101101011111110000000110101001011100011000100000100110000111000000100110001110100101101110101001110111010000011010110; 
out3543 = 128'b00110101000000110001011111110001000000110101010011110101110100011010101011010001001110101000100101011001101110011011001100100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3543[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3543, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111000011000100110000010010011110000001000000110100001000001100000111001001101111000111000001111110000111101100000001100100; 
out3544 = 128'b01010011100011100111100011001011110011110011110000101011001010110001000001010111100010000010101000000101110001111110111101011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3544[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3544, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110100000100100110010110011000110100001111111001010000011111010010000100100100001110011000000011000101110011011011110011101; 
out3545 = 128'b00100100100010110101010001111000110110110011001111011000101110011010000100111101010110010011011100010001110110001101100001111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3545[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3545, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110101000101100110011010010011110110101001100110010001001011000110101000001000111010111001111011111100111010011010001001100; 
out3546 = 128'b10010111110101001110000011110110001011010111101001111111110111010011011101100010011000101110101101100101110011000100000010011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3546[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3546, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110010010100010001100011111010001000001011000111001110011100101101011100010011111111001100011111011010000010101010111100101; 
out3547 = 128'b01010110111000101110111000100100110100101010110100010111001011000101111110010111111010001001100000000101000010111100101010000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3547[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3547, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001111001010100100111000000001101110011001101000001001001111000100100010111100110100000011001100001111001101011011010001011; 
out3548 = 128'b00000000100011100010110110011110101000100100111101100010110010010111111011101010011000100110010101010010000011000111100000000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3548[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3548, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000111110110110000100111100001000110001010100111101011100110111101111011000110000100011000101001011111110001110000111010111011; 
out3549 = 128'b10111111111111111000100000010101001100001100010111011010001010011111101000110110000100010001100101001000000101000111100111000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3549[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3549, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001001111000001100011011010001011101010101110100100100001100011110000100110110001110100101001001000101001000110011101000001; 
out3550 = 128'b00000000011100110001110011101000001011001001101100000101010101001110100000100100100000110100010000111100001100011100010000111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3550[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3550, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111111101011110011101111101000111111100000111000010000000100011011100101000100101000000010010111000110010010110000100001001; 
out3551 = 128'b11011011010001011111000011000101110011101110011010110001010111100010011101101101010101001011011101001100001110000011011011000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3551[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3551, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011000001001111010111110111001101100010000010111111011001100010101111000010001000010011111100010001100010010010001011100000; 
out3552 = 128'b11101000011010011100111010100001010010111000001010110000000101101101010000110101101001011001010101101000011011101110001110000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3552[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3552, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111111100101001111000100001100101010111110101001101101001001001110001001100000101111011101111001010100110110011011011010100; 
out3553 = 128'b00100100101001110000110110000001111000001000011101100100101011000000100001001000100100011000000101110101110001111011010011011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3553[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3553, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111010010110111101110110100111101110100001110111110001101100001110110001011100000111011110000011011011110000110011001100110; 
out3554 = 128'b11110011100111001000010100001111110001101000010111011100000010000010010000101110011101111101011011110010011101100000101100001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3554[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3554, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010110001110000110101010100011000011110010001010110101000011110111111010001110001111111010001101011101000001101111110011100; 
out3555 = 128'b10110010001101001110111110010001011010000000110101011111010010000101011001111110101001010001101001111101111001010001011010011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3555[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3555, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001101010101010011010100100000101010110101000110100110100010100100001010110100101001000010000011011001010111111001011110001110; 
out3556 = 128'b00010001101111011010001111101000101111000101000101000000001000111101011001100000011111011100101010110011100101000110000001100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3556[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3556, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001011111101100001111111000001011111100100001101001011111110011101000110100100011001111100100000110011110111110110010010101; 
out3557 = 128'b10100010111011110101001001100101110101110000010111101101100011000001010101011111101101001000010110111101101001000110000000010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3557[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3557, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110110111111111010001101001100111010011101010100100000111011101101001110101101001111101001110000100111100010101011110111100; 
out3558 = 128'b11110010011110001111111100000001100100011010000100001010011001010101001111000110110000010001110000001011110010011011101000010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3558[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3558, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100111101100110110000111001111010101000000100001100110010011010101000110101011110111110011010100001111000101110001100010100; 
out3559 = 128'b00110011100100101100110010001100000011011010000101111000101110011100011110110100110111001010011001010001101111100001001010100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3559[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3559, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000110001110010100011011001001101000110100111101011000100110101001001111100101110110111011110100100010011110001000110100111; 
out3560 = 128'b10101000101100000101000011101011110011100110010101000101111001010111000100100111101010101001000111011000100010100000001110001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3560[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3560, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110000100110000101101111100110101110100110011011110010010110100101100111000100010000100101001100101101001101111100100011011; 
out3561 = 128'b11111111000101111100011010010000111001001010111001001101110110110001001110100011111000110000100101011010101111101110110011100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3561[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3561, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111111001111110111111001100101010101000011100100110100010010110010000111000111100100101001011011110100111011110100010101110; 
out3562 = 128'b11101001001110011010111010010111001100111010110101010111001100011110110001011010100100010000111001011111000101111111110001001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3562[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3562, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000111111100001000111100011010101101101000000010010011111011100010101101101101110011011111011001100000011010001111110000111101; 
out3563 = 128'b01111100011000000100101111110011110011111010011001111111110000100110001111110111011010011010100110101000110110000111001111011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3563[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3563, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001001001000100100100110110111011010011101111001000000111011101010000000011010100001111000011110100010111100000111010010000; 
out3564 = 128'b01111010101001011011111000101111000001111101110010011111101110100001101011000111001000111010111011110000000011000001110011100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3564[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3564, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110010011011100101000100010110001001000111000010111000101110110101101110110010001111001101100100000010100010000101000101100; 
out3565 = 128'b10000010010001100011110111000001000001011101100011111010000101111101100000111000010001001100111011010111110110101011011000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3565[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3565, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010110011110000011100000001001100011001000111001111101010111100011111001110000001111101101111111011111011000001011111001011011; 
out3566 = 128'b10110001100110010101010010011000011100011100100110000000011010000011011111010001111110011111101001110101111101000010110000101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3566[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3566, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001010000001100111101000010100101101011101000111111100110101010000001110110001001001000001001010010000110000100011010000110; 
out3567 = 128'b11000010110010000000001010011101011111010100101111011010111010101001001010110010111001010101001010001101110100110100100010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3567[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3567, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100100011101000011011000010011110111110110011011000010011111010111110010001111110001110110011110100001011011100101000000101; 
out3568 = 128'b01100100000100001110110110010000101100101111111101010100110100010001000110011010111000100100000110010110101111100100011111111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3568[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3568, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001100110101100110111001000010011000010101110001010110000000000011001001100101111110100111001100100000011001000000000000110; 
out3569 = 128'b10101110010110010010011111000111100001010111001000000111001011010001010100110110101010010010101011001000010101010001010101101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3569[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3569, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011001110001010011100011100110110110000000100000110110011101111110100100011001000001010000010101010010101101000011011001011110; 
out3570 = 128'b00110000000001101000101010000010101011010101000110100011011101100001011101001000100001011101010000000010000001101001100000110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3570[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3570, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101100001110001101000101000001110011011011100011100110000011111110101000000000101000101001110110011000000101001010101100100; 
out3571 = 128'b10101101011101000111001010101010101011110111111011110110110110001011011101101100101001110010101010101010101100000011011011000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3571[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3571, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111111010101001010010110110011000010010000111011001101001000010100111111101100011011000000111011000000011010110010011111001; 
out3572 = 128'b01111100101100000011000001000100000111101010001001011000000011001010110011001101001001110100001011111001111110100001001001000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3572[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3572, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111100110111100001011000100111101001011110011101010011010010100010110010001011111010001000010000011110011000111100011101100; 
out3573 = 128'b00001110110110110010011100101110000100100100000011011101111100110010001111001100010101111110000000111001001000010101000000001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3573[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3573, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100100110111001010011100111101010111001000010101101100010100011101011101100101110101111001011100001011001001100011100111100; 
out3574 = 128'b10100111011100010111001001111111100001011110101100011110100111011011110110010110010111111101110000001100010011010101011000000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3574[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3574, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101100011110110100010101100000010001010001010111010010101110111111000000000011010010001110001001110010111111010100010000111; 
out3575 = 128'b00100000110101100011011001101110101111001101101111101000100101010010000101000011111111010001110110100011111110010010101101001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3575[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3575, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110110010110001000001101010111101000000010100101000101101100011000000011100010000000100010010011110101111011001010110110011; 
out3576 = 128'b00000101011110010010100011110001100100000110100000001100000000010001000100111000011101100011001011011001000111010110001001010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3576[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3576, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001111110010110111110100000111001101001110011110001000000001101010101001000101001000111100111111000000001010110111001011001; 
out3577 = 128'b00110011001000000010100111111001010111110100010010111111010110001110100101110111010010000100010111000001001011100111011110101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3577[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3577, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100111010010100001010101010100111010111111011110101100100001011010010110100110001111100100101000101011001100010111001010110; 
out3578 = 128'b11000010110010101010001110011100101001101000110110100101000100010000010101100001111111011001010001110001011001010110101101110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3578[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3578, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001000011100011011001000101001101101010010011100101111101011110110101100110100011111001101101000011101100001011001110101010; 
out3579 = 128'b10111001110010010001000011000011001101010111110100001101100101001001111000101000011010111111101000111000101010010110010101110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3579[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3579, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001000111010101101000000101100001100000000010001100101000110011011011010110101011011001010101000110100000010010000001100110; 
out3580 = 128'b01101010010100011000111001111000000101110110101101101101110011010111011010110110000011010000101011001000010001001100001001001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3580[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3580, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011011110010000100011111011101001010111110110001011101111100001001000011000000001110011000111110000011000111000100000101001; 
out3581 = 128'b01000100011111000001001001011101000010101110010001111011010101001010010110000101110011010010101011000111011000100011101101110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3581[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3581, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111100110010000100101000000000010001010010010111001101101100111100011101011100101111000010001011001010011010001000110101000; 
out3582 = 128'b11111011100001101110101110000111011011001001011011111001110111110001000010010011110101010100011011000000101101001001100100111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3582[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3582, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110110100001001001101011011000111011100010111111000010110111001001101100000110001011011100000010111111001011011100100001010; 
out3583 = 128'b10101111111110011111101101000110011010111010010011111001010001100100010001001010000100011011001000011100111001011100001110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3583[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3583, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000010100100111011001000111001100001001001001010011100101101010111110010101000110111100000100111111101001110101010011100000110; 
out3584 = 128'b10001101110110011100000010110001100001110100010111001001000011100011111111111001100100111111000111100110101010100011100001000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3584[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3584, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000110111110010000010100111011011001010000001101001001010111111100011011011101110011000011010110111011110110101110010000101; 
out3585 = 128'b01010010100000010101010011110111010010111101100100110111110000011000110011110110010010110010010011100111111000110001100010111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3585[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3585, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000010010100011001101100100010101011111011111101010101100110011100001100000011010111001011000110101110100101101001111100010; 
out3586 = 128'b11011011100001110000001100011110110111100011100110001001000100110001110100010000001001111101011100100111011010100110100101011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3586[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3586, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010000001101111101101101001001010111010110001010110000111011110100000110001001100100000011111100010010000100100111010001110; 
out3587 = 128'b01001011110111011100101111111011011010100111010010001110101110111100110011101011101010110101001010101110100110111001110101011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3587[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3587, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011010001010010101100100100101111110000001110110000101000001101010110100111110101010111100010000110011000000011001101000110; 
out3588 = 128'b01001001011110010101111001111000011111001000010011101100011000100010111111001001111110011111100011000101100100001001100011001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3588[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3588, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001110110000101100000000010001111100100101000010100101001001010001001011001100100110100001000011000001110010010101000110001; 
out3589 = 128'b10000101111011000001101000101010100000001000001011011110110001000100010100110000101010110011001101110111101101100100110011010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3589[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3589, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100110011000001110101111111010100111010011000000000100110001000111100100111011111010000101011111010000011110001011011110111; 
out3590 = 128'b10100010001000111110100101001111101101101001001100010011000100011101100011110011011000000000011100101011011011010101011010000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3590[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3590, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111111101010101011101110011100011101010111110001111010111010101010110011100000010010111110001110110010001110101101000001100; 
out3591 = 128'b01110101001110110101101010000100110011000001111000111101011111111001010101111011111000101101110110011001110100000100100101010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3591[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3591, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101010110101110001111000110111000011101110000111011101001001010011111011000111110100000010100000001101000000101011011100011; 
out3592 = 128'b11001110010110110000000110011101001101010110111010001001000000111011110110000100000011011100110101001010010111111101100010001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3592[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3592, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100101010111101101111100110001000110010101100110010000011000100000110111101000010000001110001010110010001000000100101110110; 
out3593 = 128'b01101111111000100110000000101010001110101101011010011000111001111011001110001001000011000100001000100110110111111011000001000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3593[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3593, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011100010110101010000001100000011110100101110010000000100111110101001100010100100000111000000100001000011100000111000010101; 
out3594 = 128'b01100011110101010010101100010110010100010001010001101100000001101000001000111001110001111100001000111011011100010011010100111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3594[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3594, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111100100111111101011110100010000010000110101011101001111111011000010011000100111000011100100101001001111110011010010000000; 
out3595 = 128'b01100111010011100111011101010101110000011111100000010110101110111101001010111010101100010110111011111010010001100000100100000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3595[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3595, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011101101110100011010100001111101011000110110010000010110011011111001010011101111000011101101100111001111000111110010011000100; 
out3596 = 128'b00111010111011010101101000000000111101011010011000100010010101000011101110011010011100111011011101110111010110001001110110001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3596[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3596, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100000000101100101110100010011111010101101011110011010001111000000101001001000111110100101111010100011011111000010001110101111; 
out3597 = 128'b01100001100101111001101010111100010000101001101001100101011000111000101100011010100110111101000000110010110110111011100010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3597[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3597, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101010010101110101110011111011011100000000001000010011011010110000001010001001000110100011010001101011100001011000101000001; 
out3598 = 128'b01101111001101101010101010011011101111000101010011110101000110000001000111111101101100010000100010101111001011000110000011000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3598[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3598, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100011001110101110110011011000011110110110001101011110011111011110101010110001100001000011100000000000000100100001000011110; 
out3599 = 128'b11100101111011101100001101111101011011010010000110110010010110111011010100101000001010111001101110000101011001001100010010011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3599[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3599, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101000011111100110101011110101000000111111110111111101110010101011110100111100000100101000101100011110111010100101000000010; 
out3600 = 128'b01111000101111110001010111010100010001111100101100010011100110001011001111101010101110111100101101100101110001111011001111101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3600[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3600, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000010111100010010001001101001110001111001011000110111011000110101101111010000010111000100101010000100110010111011101110010; 
out3601 = 128'b01000111010001000111111101110000111000011110101001001011011101111110110010000101111011111111001011001111100110010010010111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3601[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3601, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110011011111110011110101010110010000101101000010011110001101101010000000000011000011111110000110111011111010110111000111001; 
out3602 = 128'b11000100101100001010101111000000011100000100010110111110101100010111011110111101001100010010010101101001100010100000100110011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3602[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3602, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110010000111111001001110010011011111110100001111111000100010001110111110110001111000000011101110110001101011111101011000101; 
out3603 = 128'b01010111001010000101000001110011001000111111000111010010101101010100001111111010011110011011100001000011111000101000000011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3603[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3603, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011010010110011010101100010101100110011110001100101101010010101111100001111011111101110100110101000001000001010010001100111; 
out3604 = 128'b01110010111111000100100001001010100101010011111100001110101010110101000111111110010100000001010111111010100101000110010111101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3604[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3604, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010100010110101100110110010001100110010110001101000100000011001110100001001100111111001000001101000001001101111110100001111; 
out3605 = 128'b01001101001101001110000101100101001001111101010001000111001001001110111011010001111101001110111000001000001110110011001001100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3605[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3605, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001100110111011000000100001010111110001110100010000110100000110100110101111111100111010110111111111111011000000010100001101; 
out3606 = 128'b01111000101011011001100000001011110110101010000000111011101010001111111100100100100000010101001011100000100100010110000010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3606[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3606, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101100101010010110110110010111101101101100111011000001010010001001111000011000110001011100111100101001111101000110000010011; 
out3607 = 128'b10010010010000011000011011010111000011110001010001000001110100101111101100010001001010001101100101001101000010010100001010001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3607[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3607, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100101010001001010011010101001000011000110011101110001011001011011011111110100010000101101001100000001100010111000111111110; 
out3608 = 128'b11110010111100001001011011110011000000011100101000000011000000101001110011111011001111110011010111101001000111101000101110110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3608[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3608, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011001111000111011010111100100101100101111111100100110001101000100011010000111101011000111000010101011001011000100100001101000; 
out3609 = 128'b10011100000010010010010010001100101111100100110110110000000011000111101000100000101011100111110101010110100101100000100011110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3609[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3609, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101011010000001110010110111101010101000000110111100110011100101100011101111100011000101110000110010101010001100010110010000; 
out3610 = 128'b11101001100111101101101010010010111001101011110001010100101000100001110000111000100010001011101100001110000011001000100011010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3610[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3610, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101101000110101101110110000011001101110001101101001111100111011001010100011111010101011111101011111111011001000100110000111; 
out3611 = 128'b11111101001010001000001111110010000000100111000010011001111111001011101011001000010001110101001100011100001100000111011111001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3611[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3611, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011101100110110011111111100010110011110001110111101010011100100011010010110001101101001001111010000011100000011001001000010; 
out3612 = 128'b01001111101001010001011111111100011000001000000111000010111101101001011110011110000011000010001010001000101101011010001001110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3612[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3612, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001110110110001011001001101111100100101100010111000010001000100000011100000110000010011101001010110010010000100000000000110; 
out3613 = 128'b00001000010100110001101100111100011011110110011000101111111010111101001000110110100011011000100100010010111000100110010110001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3613[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3613, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000100100111011110101101110000110100101111010010100100110111010000011110001010101000110111111011000001001111100000111001010100; 
out3614 = 128'b01100110111011000111011101101100010010100000111011100010110101101000000101101001110000001101100111000001001110100111000010110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3614[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3614, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001001011000110001010100111110000101100010111100010100010010010001100000111111001011010000011101100011001010010001101101100000; 
out3615 = 128'b10100011001110010000010111000011101110100111111010111010010011111011111100111011000000101110001110011001100111110100011101101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3615[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3615, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000101001000111100110001010000000111001101100110000111101101111111100101101100011000011100010000000011001111110001010001111; 
out3616 = 128'b11110101111001011001110000011011001100010101010101010001000110010000011000111011100011101001011001111100011100111011011000011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3616[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3616, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101110011011011100001100011111011001000100110101001111100001110100101001010000111011011010111001100010100001111110010000000; 
out3617 = 128'b01101010010001000011100011111001100010111101010111110100000100101011000101100110111011000110110000110010111110000001111001001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3617[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3617, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111100010010001011110010001110101100010101111001111111101000101100001101101001011011010100111111010001000000000000101111110; 
out3618 = 128'b11111100100000111011001010110010100010100001100100110100000000100100101111101000010110000000010100000011110010101100100000011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3618[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3618, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110111100001010011010000000011111111100110110011110001000101011111100000101110000010111011010001100001100111101110000011011; 
out3619 = 128'b11101000101111100010010001000010010110000000011110100101111110000011111001111000000100011000000100100101100011100000010110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3619[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3619, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001111011011011100100101011000100001101000110011010101111100100001000001100110001110011110101000111100111110110000000001000; 
out3620 = 128'b10001000001110111010010111100111111001110010111001000001100011100011010011100111011011001101101011010001011110110110111101100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3620[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3620, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010101110010110000101101011100011101101110010101010110100100011111110011101111001100001011011001111101111011000011011100000; 
out3621 = 128'b01111101110110100011101001100010111111001001111111100101000011010111101100011100101110011011110110010101011011010001110111100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3621[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3621, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101100001100011010101001010000100111101111101111001100001000000001001111101110000001111001010111111000111101000010110011001; 
out3622 = 128'b00110100000010100100110110001011000011011100010101010001001001110110101010110111011111100010101010011010110110000001100001111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3622[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3622, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110010011010111001100001001110011100110110110110110011110100000001100110011001111100101011110110110000010111111001011000001; 
out3623 = 128'b10110011001001100110000110000111111010001101100110111100011001111101100001011010000011110110000100100111101101100100101010110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3623[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3623, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101111000001111100011001011110000011101010100110110010110111000101110110101111110100111111000001010000011001011111010101101; 
out3624 = 128'b11011111100110110111001100000001001011011110010100110000110001100001010011110010111010111000000001010110011100001111001000111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3624[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3624, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000000001110010111110111000010110100111110100111110011000000001001010110001011100110011011001010101001100000111000101010001; 
out3625 = 128'b11110011010111110001010101011001111001001011111110001000110100001100011001100110110101100011010010101001011110111000111011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3625[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3625, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000011110011000010100111000100011001010011101011110010001000111001010110101100011001011000001111001101011101100101000100011101; 
out3626 = 128'b00111101010010011101000101010100011010110010100011101001101101000011001111011110011001010111101101011100011011110100100000110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3626[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3626, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011101110101111010001110110010100101011101010110001110110010001101101100110001100101001001101111011001100010000111011100100100; 
out3627 = 128'b00101000001001001001001111001011101000000011011100000001000101010111010111110111111101111001011110010001111001110101111111100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3627[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3627, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001110111110111110101001101011100010011111101001010011111001110110110100011101010011000100011111000110010100101101101101011; 
out3628 = 128'b11001000111000100011000000000110011101011010000011110000100001111000110110101101110111001011001100110100110001100111111011011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3628[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3628, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100000111001011110000100011010100111010111110110110101100011000101000001101010101110011000011101001010110010010111001001010; 
out3629 = 128'b00111100110001001001111000100000100000011111001011110011000110000010100011010101011110101001011110101100111111111000000110011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3629[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3629, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011010100110001000010110010110101000111011001111100100101010100011100101010111001010101110011100110110111001101010001111011; 
out3630 = 128'b11010101000100001101011111100101010101011000001000011110001110010010010100101011010011110011001101000100110101011000010001100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3630[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3630, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010101010000100000110110100010110111101010100110111010000001101100100010111110101011011001001001001011101100000101100000101; 
out3631 = 128'b10001010100011100001000101101101001101011100001001101010110100110001100111101010010110110111101101110001000101111001100111100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3631[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3631, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111111001001010001010010101100101001010100101010101010010011010011101011111100111111011010101110101001110101011001100111010; 
out3632 = 128'b00101011110011100001100001111011101000111111011001100010101010110111110101110000000111010101000000011011000001110001100111011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3632[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3632, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010000000111100111111000001011101001100101000001110110001110100111000001100111010000110101100100000000010111111101101000001; 
out3633 = 128'b01000110111000110111100010110001101010101010001010100011001100110011011111101001011000100001111100010110110100000110110001100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3633[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3633, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100100111100101011101011010110110111000101111011100110000100101111010110010100100000011000111000111001010010101111101110100; 
out3634 = 128'b00100001011110010110011000001010100000111001100010100001011111101111111001000001100100000100110011101111101001111111100110111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3634[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3634, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110110100001010011101010110001111010001101001001111110111001010111100000101111011011110010010101101000010011001011101100101; 
out3635 = 128'b01011000000101010011010111101111001100010011101101111001000011100100110011101011000001110000111101011101101011010010100111100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3635[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3635, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011100000100111011101011001110111000110111000101000110101011010111001010100111110101101010101001001011001101001011010100001; 
out3636 = 128'b10101011110110010000001011111101010000111100111000011100110001011110001101110011110101011011100000111000001010010101101001010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3636[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3636, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110110000010010111001000010000110011010000100010110110101101111101000110100000001101110100001100111001011000110010100111010; 
out3637 = 128'b11001100111111001110010110000000101100101001000111001001001101001100100010110010100100011101111001000101111011111111110011011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3637[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3637, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111000011010000100111100110101101001101111110100110111010100101110010011111101001000000111010001101001011100000100100001111; 
out3638 = 128'b01000010001100011001110010011000011010011011110001101101001011110101011000101100001010100100011110111110100111010101110000001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3638[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3638, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001001010110111101000101000110010111100110111001000000100111111110010100100010011001011010110101111011110000011101000101110; 
out3639 = 128'b11111110010010011100000000000010111010111100001011100101101101001101011111100010111010001011001011011010010011011010001000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3639[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3639, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110100101101100010101011111011001010101110101110000000000010000011100100111011110111011110011001000111111010100001100000111; 
out3640 = 128'b10010001101001111001000111110010011010110111100000011100111100000011001101100010000110110001101000010111101001100111101010101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3640[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3640, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000111001101101001110110110100110101000100101011111111000000011100000000011111001010111000001110010110011010101101110101100; 
out3641 = 128'b01111010010001010100100000111111101001100110100010111101100100101101011011100100000111101011101111110100110011111101010011111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3641[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3641, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101001001100001011010110001011111010001100010011010110001011110011101100001010111111001010110001100010001101010011001110111; 
out3642 = 128'b10011010011110110101101010100111001000011000001100110010101100000101101110100010111110100000011111010100101101001011101110000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3642[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3642, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111010010111101010100011100101010111001001111000111000101001001100111001011110001110101101100000011011110001011111101111000; 
out3643 = 128'b11010010000111000010111100111101101101111010111101111100010010001000101010100100111100100110111011110111010010010100110110101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3643[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3643, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110011111100011111001000001101000111100101010111110111100110001011111101011001011000000110010000000111001001000011111111001111; 
out3644 = 128'b01000001110011101010010001000100001110010001111101101111100010110001000001001101111111101100101111100000111000000101111010010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3644[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3644, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011101101100000100100111011001111010010111111100000111111001111100001001001101001011000110100111000000001111101001111011111010; 
out3645 = 128'b01110000010011100110010001010100111001111000000111011000011100000010100111100010010000101011110100010111111000000011011011111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3645[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3645, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000001101100111001111011100100110111101010001110001011100010001010100111110011000010110010000111111000010101000000000010011; 
out3646 = 128'b00110101011101111000101001010100000110001001010011011110100000111000000100001111110001010011000010101100011100000111110100011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3646[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3646, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100110010101010010110011111011111011101000011110001000010001010100101011010111011001001010001100100010011101100111001011000; 
out3647 = 128'b01111100010101111011011101111010001100001100110011100011001110000111001110100010001110111000111001100100011100000011101111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3647[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3647, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101111010110100010001100111000100000011100111100100111011110010010110001100001110110110100101111101010110100011100101010001; 
out3648 = 128'b00100111111011000010011101011000111000000011111010000011110111101110011010100100001100010100011010111010100110001111010000100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3648[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3648, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011011010100111101111110011000000111000000011111010101101011011011011001000011010101110110001000001010100011111111100000111; 
out3649 = 128'b11110111110010010010111110011011000010111100001101011011110100011011111001011000110010101001100001011011110010110010110001111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3649[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3649, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110000111101011110000011110010011100010100001110101111100111111111101111011101011001100001111110110010110000011111010101001100; 
out3650 = 128'b10010000110101111000011110101010111011010101111010100011110001001101100110111100010010111011011010010111010010011010111111000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3650[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3650, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111101101111011000011110101001010100011100010110101001101001100011011100110000011011001001110100010010000110100110011110000; 
out3651 = 128'b10100010010110101000001100011001011011101010100010100001010010100101001000110111110111011111111111011001001010111110011100001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3651[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3651, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100100011010101101111001101010010011000101001100101101101001000101001011111000010111001100000000101110111011110000011011111; 
out3652 = 128'b11001011010010101110110001000010100001010110110001100011001011111011001010101011001000110100101111000100101100111110100111110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3652[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3652, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101110011100111001001100011111101010111110110111111001001111101111000101111011100100111111110001000010101011100011111101011; 
out3653 = 128'b01110111001000011010010010001100000010100011111111010101100011110000010001100110111010110101010011011001010010111011100011011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3653[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3653, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000100000000110010010001111111000001100010101100001111000111110101100001000111001101110111001101101000011111100110000000110; 
out3654 = 128'b10100011100001001011001110010010111110100110111010110000011001000100010010000000110110010110011101110000111011111110111000001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3654[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3654, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110101101001001001000111111000010000100000111110100110100100101010111010110101101011001110100111000001010101001111100101100; 
out3655 = 128'b01001000100100011111010001100001000010111101110001110110101111010000100000001101011001111001010111011000110101001111100010001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3655[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3655, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100000101110110010101101000001010111010100111111101101010111010010011100001100000010110101110110100010001011011001000010110; 
out3656 = 128'b00100100000000111001101111001110100011100010000101001001010110101110000011011100001010010100000010011011011110011001110111100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3656[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3656, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001100101001000110010000001010010001100100110011110010100100101110110110000010111110101111100111100100100110101010110100111; 
out3657 = 128'b00010001101011110001100111010001111011111100010000100100010100111101010100100100101001101111000101010110001100001010010101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3657[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3657, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001010100110010101111101100111010100011101101000000010011100001010101000111111111100010110110101010010110110111011111011101; 
out3658 = 128'b01011111110000000110100110010010001110111101001010110001000110011010101101111101001101101001100000001001100011101001010001100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3658[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3658, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000001111111101111110110101010010011100000100110001110010111011000010101010101001000010101101010010100111100101000111001111000; 
out3659 = 128'b11111010111010011011101101110101111001011101010000101010110011010000111101010010000000010110111001111011000000001110100100100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3659[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3659, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000010110010011000110110001010000101011111111111101111101001010001111000111110101001101001011101001011001010011000100110111; 
out3660 = 128'b01110111011011010011100111001100010100010010100101000101101110111000100110011110001111100001000011011000111000100000111001011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3660[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3660, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001111100101110101111011010011011011111101111100001100000110001110011110110010101111101111010011011011001010000000011000001; 
out3661 = 128'b00001100110110111101001000010111001100101101000111110001111110110110011001010110000110011110100100011110100000101001011001001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3661[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3661, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000011000110010001100101000001000010011011111010111001100100011101001010000011000111110110111101100101011010111101011011010; 
out3662 = 128'b00101011000000011010101000010011110000100110011001100010100000000110010101010000011110101101110101111111110100000111111110100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3662[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3662, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101111101111110011110100001101000101010101001011110110001010111111000011001100111000101100100010011111010100010000000010011; 
out3663 = 128'b10011010011010011010101010100010110010111010100001010000010010111100111010111011000000100101001011101000010100000101111000010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3663[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3663, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100100001101011110110011100100000010110011011000001111101010100101101010001000000101101101111010010010111000011001000101100; 
out3664 = 128'b01100100111100101111011001000110101001001010110010101001101110010001011100101111011000010010010000000000001110000100011000111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3664[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3664, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111001100101011111011100101110001000011101010000011001001111010100011000011010000000100011011011111001111010111100000110101011; 
out3665 = 128'b01110010100101011011111010010100001110001011010101111111111001111001100001101001011010110000011100011001001000101001101111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3665[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3665, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011010001011101110001011101111010011100101010100110001111101101110101111100100100010111100000011110010101100100011100010001; 
out3666 = 128'b01010010101011101011011111000001010110110011010110001011100100100000111011011111110101011011111010100010011101001010010110001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3666[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3666, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101011110100011010001101001111100101011100000000001000001000111001011010100001111101101001000110010011110000011010100001101; 
out3667 = 128'b01101101010100011101111010100111101100011110010111100111001111001111101010101011001101101001111001101001001000110000010001001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3667[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3667, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100010111110000111010000011000001100100101001110110000000111001010010001101000101100110010100001010110011010011011110011001; 
out3668 = 128'b01100110000011011100000010110101010000010110100000011111101010110111111001101001111000110101010000111011110111100011111011001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3668[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3668, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000010000000100011110100111110001011111111110001100110010001101110101110010111111101011101101111010111110110101000111010100; 
out3669 = 128'b00101010110001000110000101000100000000001011011100010010100101001000001010001111000101000110011011001010100110011000000010110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3669[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3669, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010001010101001000001110011000100101100001010001010010101010110111010001010110111010011011110001010010010100010001100000011011; 
out3670 = 128'b10100010110001100001110001000111001111110110011001010011011110011111110010100011111111101101101100001011111011111110100111110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3670[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3670, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110000110000100100100100101001000111011010100010101010101110000101110101110011110100101101001100101111001010000110101011111; 
out3671 = 128'b10010001101111000100110000000010010110000100000101001010110001001011110110111101011101011011010001101101010111001011011011000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3671[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3671, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010111101111011000111010011011000101001101011110010110100101110011111101000100111101100001001110110011011000000011101010010; 
out3672 = 128'b11000100100100111111111100010111001110111000100101100010110010010111001100100100011001110110010010100110001110011011101001100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3672[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3672, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001110110010010001011110011011101111111001111011111001010000010001100011111000100011100100101110000010001000110101001000111; 
out3673 = 128'b00011110011110110010001000000001100001110110111110001110101000101111001000110100011101011110001001010001001000001110000011011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3673[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3673, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100000010000011011000100101111111011100011001100110010011001110111110101000001001101101001110100100110010110101110101101011; 
out3674 = 128'b11111110111001001110010000001000110001110010100101000000000011010101101011110011100010101110100101101110100111111001000100011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3674[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3674, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100110001101000100110000101001110111011001110001100111001100000100010111010010001000110101011111111111010010100110011011101; 
out3675 = 128'b01111100111010001111011111100001001010111110001100010011101000011101100011001000001111000100010010110001111110001011000011100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3675[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3675, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110110010100111001101100110011001011111000111100101000100111100001100100001011110101111010011001110110011000010101110001100; 
out3676 = 128'b00011110111101101110111110101100111010011101111010001100011010111001001100110111000110001000011101101011010000101001101010010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3676[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3676, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010001110111111011101111111001100110011111111010001100101011110011100111111010101011011001111010000010010110010010001010111; 
out3677 = 128'b10000011010000101111011000110010011001000100100101011111011011100001111010010001110111011001110000110001101011100001100001000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3677[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3677, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100001011000101111111101101100001100010011011010100111110010101010010100100101100110000010011101010011100101101011110010111100; 
out3678 = 128'b10110111011000111001001110010101111111000111111010011101101111100101101011001011010011010001010000000000110111110000101111000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3678[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3678, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001110100000010111101001101100011111100110110011110101010100110110000001000101100111011110000001110011011000000100110110000; 
out3679 = 128'b01101110101100100000110001011001010110110000101000010110000011111101110001011101111101010110011110111110000111100010101111000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3679[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3679, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100111100000110011100110010000001011100000011011001100011100000110110011001111100010000110101111011010011111011101000011011; 
out3680 = 128'b01011010011100101010100011100111000110000000110101010010000000000010100000000100010100110001111011110001011101111010001010110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3680[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3680, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101101000100011010101100000001100000110110110101010100010011000010000101000010100111111011110001110001110100111000001011111; 
out3681 = 128'b10001101110111000000010001101011010111001000000001111001111010010011001001000010111000010100100001010101010010101110101010000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3681[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3681, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000100111111111110101001110110100001010111011011101000100010100100001010011110011110000011001111101110101011101000110110101; 
out3682 = 128'b01000010101110001010000100101101001101000010100011101110011011000010000110111110001111111010011001100000000000010000000110000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3682[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3682, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001000101101101001110001011010001111010110111110000111001011111010001110001000001111010100110110101001010110111000010110101011; 
out3683 = 128'b11011000001011001010100110110100111010001100101100001111111010000100110010110111101000011010011110001110010110000001101000000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3683[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3683, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011011101111111100000001000000001011001000100011110011011001000111010100110011000100111010010111101001100111000100101101110; 
out3684 = 128'b01001111110000010000011011100100100100001001001111001111101011001011010000010111010010001100110010111001110001110100000011001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3684[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3684, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001110001011110010001101000001011111010010110110101101011111001001010100111110001110111000100000100001000110111111101111100; 
out3685 = 128'b00001111000101010110110001011001101000010110111111000001110100110000111000100010011111011100100100001100001000110001011001111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3685[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3685, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010010100101100011101010010011101101110100010001101101110001101101111111111001010000010000100001000101110010111101010001101111; 
out3686 = 128'b01111100010111011011101111000000001101000001011001101101011110111101100010011001100101110000110101100001110011010001111100101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3686[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3686, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100100110011010001111101110111001100111111100001101110111110001111110101100111101101010111100110101110110100110011010101001; 
out3687 = 128'b11111111110100111011001000101000100001011110000010100010011010011001000010111100010110010010110111011110110110101110111100011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3687[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3687, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011101110011011011011111111110110110110110000100001101101011110000011101001111010111000110001000011011011111111010001000110; 
out3688 = 128'b11010110100010001000001100000001111111010011001110101000110011001010010000111000000000101011111110001011101110110100110111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3688[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3688, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101000001000011000001001001111110011000000011111110000111001110010111110110000010100011011011010000010110100011100110011111; 
out3689 = 128'b00000110010011110100011010101010000011100011000111010100100110101011110111100011001100111000111110100010100110011101011001101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3689[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3689, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011111000100010101110001001101101111111001010100011011110111010110001000001011101110110010010111111011010101101111000111010; 
out3690 = 128'b00101011101000010111111001011100011111011110000110100011001101000111000010010101111110001111100110011110110110000011001000001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3690[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3690, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101111111110001011101110001111010011110110001111111111100101111001101001101110100010010011010101011101110001001100101101011; 
out3691 = 128'b01100000001101100000011011111100110000101100110000011000010110011100110011011111010110101111101011101111001101010111010110000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3691[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3691, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111010000100000010101111110011000100000101010111101000011110000100000101101010010011101010100101101010101001101101101011001; 
out3692 = 128'b00110011100011110100101101100111101110000011111100001110011001101110001101011001000011110111111011101010010111010110000001010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3692[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3692, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111110111110000010011100100100111101110010111101001011101000001110110100111111000111010011001011001101000110010111011000110; 
out3693 = 128'b10111011110001111011111100101111001010110110100111010010010010001100101100111101001001101100110011000111001000000001000010100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3693[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3693, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110000111100000001001011000110000110001010110111110101000011000000011010001111110110011110101001111101001100101100001010010; 
out3694 = 128'b00001001011010001000100000000000010010100000001011110011000000111011011100000100010100100110001001010011101101100010111010111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3694[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3694, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001100010110000010010101001101011100111110100100000001111011100101101111011000110100001000100101001100000111110001100110101; 
out3695 = 128'b10110111101011001011000000111011101001111011000010010101101100011111001110100000001000000010000100011101001000110111000101101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3695[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3695, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100000101110011000110110101001000000110111001101100001100010111011010111100001110100011001011011110100101011000001100111000000; 
out3696 = 128'b11011101001100110010001101111000010001011100011010110101101001001111011011100001010011011000011110000001101011101001100000001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3696[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3696, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100001100111101100000101010110010001111010010111111100100001011100000111100010000111101100111000100101000100001110100011101110; 
out3697 = 128'b10111001000000101100001001101100100001010000111101001111000010100101001000110000100100111011100100110000111010011111001111010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3697[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3697, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111001000000010011111000010110001010010000110110011110011000100100001011001010000101111011101011101111110110100010111001111; 
out3698 = 128'b00010010011101111001001000001100001000111111110111110000111010110101011101010100110100111111011100011001101010001101100010010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3698[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3698, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110011100000101110110110011101100110101010010100010010000100111101100001111110100100001101111101001000001010100100000001101; 
out3699 = 128'b01011111101001101111111011100001101001000010101011101110011010011010000011011101100111111010001110001011101110000101001110110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3699[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3699, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111110001001001101000010001011110101110000000010011010101100100110010000000111011010110111010110111101110110011011101011100; 
out3700 = 128'b11000101010001001010011010000111011001101000000110101000000101011000110101111110110100101110110001010100100001010110011000000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3700[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3700, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000110101010000100001111000101111010010001011010001110101011110100000101001000010101001000100001101101111110000101100011101; 
out3701 = 128'b01001101011111101110111101110011000100101100010001111101111101010001110011101100110010010111001100000000101010100000001001100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3701[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3701, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111001000001111101111100010101000011011101000001111000011110000000100000100101111111010001011010000100101001100110000101110; 
out3702 = 128'b00011001111100110111010111000001001101100110000010001101101000110011111101100110000011010000101111001100000011000010001100001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3702[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3702, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001010110010111010001110010101011110100010111000100001111101001101010111000000000001110101001001110001011110110011010101001; 
out3703 = 128'b10111110111010001111110001101001100101111111010100111111111111001000111100011110000111110010111111010010001000101111110000010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3703[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3703, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101000000010111111100111101011000001101101110101010010000101111111010101111010101000011011000000011100100001000100001010111; 
out3704 = 128'b00101000100010110111000110101000111100011011110100101010011001010011001001011010110001001110110010101010010001010011101101010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3704[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3704, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110100001111101110101100011101110110001010111001000000101100110101110011101010011101110111100001001110100011100001011111101; 
out3705 = 128'b00011001001010000111001011110010010010111010000010110011000000110001100000111001100110000100111010011100100111011100001111000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3705[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3705, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100111100100110001101111000000101011101110010000110001100101111010110111101010100110101110001001011011000010011101110010110; 
out3706 = 128'b01011110110011000010010000010000101011000001111110101100000110000100111111100000100100010101000011100000000010100100011111010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3706[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3706, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000000001101010111111011010001100011100111100000101010100101100101110111101110010010001101111101011010100111101011001110001; 
out3707 = 128'b10010000110011100001000101001100110110110110111101001011100000101000111110111001011010111001000100110100011100101100011101111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3707[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3707, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100101110011111100101001110110100100101100111000001000100101111000111011100001111011011010100110010101110000110001111101100; 
out3708 = 128'b00100000101100010010101101111100100001111010010000110110001011001111011000010101010101101100111100010010101001111101011011110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3708[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3708, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110110111101000001110100111101100101100101010001001011011010001111100100000111010111110011011111101111000010111001001110101; 
out3709 = 128'b01011110011001111001010100010000001000111100110100000100000100001110111011010100111001010000011110001001110010101110010010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3709[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3709, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001101100001101111000111110110101001001011101001011001001111111110100100101010010110100111101001011110100101110010011110110; 
out3710 = 128'b01001111101011101101010001100111001110011100011100110001011011111110110010001001111011010000110110010101101100100110010111110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3710[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3710, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001111110001001010100110000001101100101111011101010101000010101000001011101011110111110001100100011100100111000011011001011001; 
out3711 = 128'b00100111001101101001000011101001000010110101110111011111001111001011111011001100111010000100010010001101100110000101101101101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3711[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3711, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110110001110101010001000100001011100000000010111001000010010011110001110001011101001110001101000100001100000110110000111100; 
out3712 = 128'b01011000111101111011110111001011000010111000010110000111111111100000101011000101100010101000010001001001011010100010001111110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3712[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3712, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100000011101010101101100011111100010000100110110101101111011000000100001111101011110010011000010011110110101001100010101101100; 
out3713 = 128'b01101101010000101110010110110001010111100100101110100000110110001100011110010000011111110110011000010011110000101101100010100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3713[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3713, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101011100010100100010011011010110101110010011101001001111101111100010101100101010110110111111001100010111000100111110110011; 
out3714 = 128'b00000100101101011001101110010111001111110011011111111010111011110010110110101111000110110111000001100110010100011111111100010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3714[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3714, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011001001011011101101010110001011001011100011110101010110110010111110100000000001111100011100111010000111001100111100010100100; 
out3715 = 128'b10111101000010101010101000001110101111111000010101000111011101011110010100011101100100011010100101111001000000101011001010011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3715[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3715, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110010110010011111111001000011100010110100010100100100011001101010000101111111010110100100101110110000010101011000100010111; 
out3716 = 128'b01100100100011111011000011001110000001110000111001010111110111111101100110101101011110100011001001101000010111100001010000010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3716[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3716, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111100011100001101001110111101000111110010011110011111001000001111010100001101011110100111010010001011010000001111100010100; 
out3717 = 128'b11101011001110011111111110010111100010101001101101001100010111001110101001111010000010011110110111100111100111001111100001110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3717[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3717, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100100100101101001110100001011001001001110010010111111011011111110100000111000011010011111010100110101000010001101000100011; 
out3718 = 128'b11110110010011011100001110010000100001000100110000110010101111111011010110110001001010101101000000100110100101011101011001010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3718[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3718, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001010001001001110010001101011101101011110010011100100100101111010111010000110010111010001011101100001011010010111001010010; 
out3719 = 128'b10000001011101011101110010100100101000100001100000111010011011100101001101111100111001111010011101000111010000011111111011101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3719[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3719, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111011101000010000000101110000011010110001010100101011101011110100111010001001011010100000000001011011100011001010110101011; 
out3720 = 128'b11011011101000101000101000110000000110101010100111000001001000100111111101011101110110111110101111100010100000111111111011100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3720[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3720, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001000100100011111101100100001111010011000101110010001101000110010111110101011111000010010001101000000101101100001010111011; 
out3721 = 128'b01000110101001101110100101001010100000100000010111100000000011110001010001110010001001110101101111001110111010011110100000010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3721[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3721, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001001001111010100010001000101101000110110101000001100011000111101101110100011101000101001100010010111000100011111110111100010; 
out3722 = 128'b11110000011101111001100100111110011100101010000111101100101011000011010010010100011111110001010110110011111001011101101011010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3722[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3722, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110001111001110111110111001111100001010101100100010001101100101000010000011001100101110111100000101101110101001100010000110100; 
out3723 = 128'b01000010010111011001101100010111100011111001001110000101101110100100001100101111111101000101000100001001110110110000111100010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3723[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3723, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011010011001001011101101101011110000101011110001110111111000110011100110110111101011011101010011011001111010101000001101001010; 
out3724 = 128'b01000100100100011101111000111111101011101001010100110011011011010000011011111011011000100100111010100011010110101000101110010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3724[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3724, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010110111100011100000111011010101001111011010101001010111001010000010011000011000001111101110011110011101101001010011100001; 
out3725 = 128'b10100001011111110011000001101010100110001001000111010110110001001010011010111001111110110010000010001101111000011010101101100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3725[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3725, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011101001010001001100010001111000000101100100000001100001001001101111010111111110100101111111000101110001011011011000111011; 
out3726 = 128'b00110100001111111000100000001101111011100110110010001110111110110000110011111011000111000000010100011100011100011010100100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3726[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3726, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100111001101010000000000011101101110101110001100011010001011101110000100011100100010001111101001001001010101111011010000101; 
out3727 = 128'b01100111111101010000110101111110100010010101010001011101001111100010010100111111100001011011110011011101101001001110010011011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3727[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3727, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100000101100011000101000010111001110111011010010101011011010010011010011011011100000101010000001111110110000110111011000001110; 
out3728 = 128'b10110111111000110000110110011001000101010001010000001100010111110111001011101011001010000010010011110100110011110101011101000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3728[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3728, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011100110011001100001100001111011000110000110011100110011000101000101110111001010100110011001111001110111010010000011011111010; 
out3729 = 128'b00000110110110000111100110001010011010101000011001100001001011101110100010101011110110000011100000101100001111011101110101100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3729[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3729, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011101100100111101110010000110111110001111011010110110001100000111101001010111001000010110111011000001001111101110011111001; 
out3730 = 128'b00011000111100010111001100110100010010010011110010000011100111000010110100001011011101111110110001010110111001010011011010110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3730[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3730, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011010000010001001101010000001001000000110000100100101010011101001110111001110101010100011001001101100001011001011000011010; 
out3731 = 128'b10001110010001110100111001001100100101011001011101101100100011100011101010001100011000110010001011101101001101010111111101101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3731[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3731, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110101111000101001001101011110101110111010001111110001001000110011010010001000000000110010011100100001011110111100101110010; 
out3732 = 128'b01011110010001110101000011000011011101100010000011011100111100101100111001100010011011011110111110000101010010110100100101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3732[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3732, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011111111111100000011111010010010111001101111000100111011111010111010011000000001000001101011110100001100110011011000011010000; 
out3733 = 128'b11100110010000110111100000000010000011011000101111111001010011001011010000100011000101110011110101100100011111111111100110100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3733[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3733, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100111110100110000111110010100110010010111000010111110010101100001011100101010110101011000100111000001011110000010101110110; 
out3734 = 128'b00001000110110010111000011010111000101000001000110101001000110101111100101110001010010110101011001110111100001100011101000010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3734[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3734, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100000001000011000111111011100101100111100010001110101011011110010001111101000111000010100111011110111000110000101111000011100; 
out3735 = 128'b01001001011000001101100100101001011001101111101000011011011101010000110100110111011100000101111001010010000011101011000000010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3735[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3735, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100111010110110001011000111101011111001010111010001001101111010101001111101010000101000011001100111011000110011010110110001; 
out3736 = 128'b00110111101011011001111011010000001001111111011111111101111000000001110111001000001010001111100100111001111101010010110011110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3736[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3736, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101111100011001011011000000110000101001010000100111000001010001000001000111110101001100011010110011001111100111110110000111; 
out3737 = 128'b01000011101010111101000011100111101100111001101011000101011111000100011111011010101000000110001100000010100110000010000011101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3737[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3737, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101110011110010101010111101110101101000101001000010001111011010101000110000100110100001101010100001010100000001111100110011; 
out3738 = 128'b11100010000101011001000111001110100001111110001111100100110111000110110000100010010101111110110001010101010101011111101111100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3738[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3738, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100111011011101110100010110111000011100000000100111111011111110001111110100100110010000100010111100001011011111000111100111; 
out3739 = 128'b10011101111100011100000011010011100100011101111111110111011010001001010100110001111001100110001111110111010011010100100011001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3739[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3739, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001010001101010000000110001110010110101111100111001101001111110011011011101010111000000010101100101000010010011000101110100; 
out3740 = 128'b10100000100011000100100000101001000000011001101010101101111010010000000000001011111001001101100101001011101110010001110001101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3740[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3740, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000010001001010010001010011010000101111010010111101110110100011100000010000101100000000110110101111111011101101001010000111; 
out3741 = 128'b00010011001111111101000110110101011001011001111000001000111101110101101100000000001001101001011111100100010100010111011000101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3741[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3741, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010010101101100100100100010101001001101101100001011110001101011001110110010111001110101110100011101010100100101110011101010100; 
out3742 = 128'b00011101101101010010010101011110011100010001111010100101101111011000111110111111101111001000001100111000010111101110111110100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3742[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3742, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110110110111110100100101111000110011110101111100110110110001110011110011110000000100011010011011110001100101101110000110000; 
out3743 = 128'b00010100001010001011001101111111001101110011100011111111000101001000100010110011010000111001101111000111001010001011000100000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3743[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3743, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011001100101001110000100011110100010001111000000010001000100110111111011110101101100111000001100011110001111111110011011001; 
out3744 = 128'b00000101101011110000101000010010100010101001110000011110011101110101110101110010011010100001000011100110010111101111111101100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3744[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3744, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100110010100100110101011000101100100101001100101011011110011100110001011001100000110010101100111101000011110110011011010011; 
out3745 = 128'b10101110111110100110000110010100100100100001011000011110011001111100100010101100011001111010010111011011000011110101101101101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3745[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3745, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010100101110111110100000000111110001011111010001100100110010010010101011000011001000110110001001101000111001100010100101000; 
out3746 = 128'b00000101011011000101111010010001100101000111011110101110000111010110001000000100010101001001000000101011010111011010010000011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3746[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3746, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110010001100001111010101010110100001001001000100101000100111110110000100100101101001100000101011100100101010111100101111011; 
out3747 = 128'b01011111100001000100011100101011101110011011001101000100000010010000011000011000000100001111100111011001000101111101111011001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3747[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3747, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110101100000010001011001101101001011110101101100000000100100111101001011100000011110011100001111110001101101110010111001010; 
out3748 = 128'b11110100101001110001010011001111011011110111011000000011111111001001010001001111001111000011011000010010011011011000111010001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3748[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3748, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101111100101011111110111001110101011010000010100111000010010110110100110000010101111100010101011011100001110000011001110100; 
out3749 = 128'b11111101010011011101101011111100100010001001100000111101100011000100101101110111101101001000011100011100110001101011011111101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3749[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3749, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001001110110000100111001110100011010110000001110011110001000100010000111011000101000100000101011011010001000101110111010101111; 
out3750 = 128'b00001001100010011010111101101011010010101011110101111000000011100001010101101000111001010010110001101100111101001001101101011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3750[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3750, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000101000111001010100110001101000010000110010011000010000000110000010000010000000000001001111111001100000111110101110101000; 
out3751 = 128'b10110110011111011011100111001101110111000110110111100101001001110111000110101101011110110111101110010010010001001010100101100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3751[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3751, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111010101010111100001110001101001101001100100000001010011110101111100000110111000101110100000110111001001111001110100111110; 
out3752 = 128'b01010000101100011101010100010010111000110111000111111000001111101000100000100111110001100011110000000010011111000110101000101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3752[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3752, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011101000011010001011011100010111000101110111001110100011011101110101010000000001010101011111101011010110010110101101110010; 
out3753 = 128'b10111011010001000111011001110101000000110000111011100111110000001101011011101000100011011100011000010000011110001100000100110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3753[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3753, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011010010010110000010110010101101101011000101100000111001011111001110001000011011101111101111101000110001111000001111101100100; 
out3754 = 128'b11001001000101100001111010000000111111110100010010001111110000001011000110110111011001000010101001010011010111100011101011001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3754[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3754, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010110101100010110010000001101111011010011100001010101000001011001010100010100001011010001001001111100101010110001111011111110; 
out3755 = 128'b01011111101100101011110100100010011100100011010100111010010010010110001111011110010011010110011110011111010011101110001011001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3755[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3755, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110010110101110011000110111101011110010101000001001010011101101011100101010101011000110010001000001101001110110011000011010; 
out3756 = 128'b11100001101110100001111110011010101011101101001111001111011110110101110011001000000010010011011110000000011111001011110101000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3756[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3756, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011100000010000000111001100110001101001101111111000111011101011011101011001100110011110001011010010000001100011100111001110; 
out3757 = 128'b11001000111110101110001100000001111101110110001010001101010000101100101100011001010001110000011110010011011000100100100000100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3757[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3757, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110110111010001100100111001010101110110001010010110110010111001100110101011001010011000000110101111111110111011110111000011; 
out3758 = 128'b01000010000101110110110110011101010100000010110100111101011101111110110101101100101000100001001010100000011001111001011110111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3758[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3758, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110011011111111110100100010011010000110101010001101110011010110111010111001010010010101110011011001111110001101111111010110; 
out3759 = 128'b10010101000000011100101110100110111110111110010001011010011110111000111001110000001100111001010100100110100001000011100100001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3759[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3759, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011010100010101110111010101010100100110100100111110001011100101100110100001110011001010110100010011101001111100100001000000; 
out3760 = 128'b00100101001000101001011010100010101010011100011001101110010100111001000110111111111011101110001110111001010110111110000000010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3760[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3760, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111110101110010010111110111100110001101110011100110001011110000101011110111111110000000110011011110101011010100001111100000; 
out3761 = 128'b10111100000001111010001111111011111110100000000010001100010010001001101111000010010011101010000011111111110100111111101010000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3761[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3761, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001101111001101011101111111011010100111101111101011011010010011000110010011101110001100010110010111101110111101011000110000; 
out3762 = 128'b10010001001001001000110111010101000110011101001010100101011100010010011010111011111000011110101100011110011000010100011100011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3762[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3762, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101001000001111101110000101001111000100100101010011111000010010110100001111101001011000110001110100111001101011010110100011; 
out3763 = 128'b11111011000101011000110000011010100100110011000011000010010101011000111110011110001000111010100111011001000011010011101000000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3763[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3763, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100010011001011011001110000011100111001010000101111101100110001010001111001010100000011100100011000111100001011101100010011; 
out3764 = 128'b00000101011001000101011100011011001110011001110001011110000111010000110000101111001100011001110111011100010100110101001111110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3764[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3764, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101110000101101110001011001010000110110000100111011011010001010100001000101101001110010010111100111001001001010101011001000; 
out3765 = 128'b10000001111011001111010100101000000011010011000110011101101011111010011011001101100010100111111101100101100111011110101000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3765[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3765, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110101001000101011111010100011011110001101010101000100011000101001000110000100000110010100011100100110000101010011010000110; 
out3766 = 128'b10100000100001010010001110100111100001101101110001100110110000011100111111001001100100010100001101010111110001110111111100010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3766[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3766, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100010111011101110111001011101101110000110001001110010101000001101001011111011101101011110000001100011001111101101111010001; 
out3767 = 128'b00011100000001000010010101100000101011111000101100011001010010101001111101001010100101010111110011111111101001001110111001100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3767[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3767, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100010001100100010001011110100001000111000101101000110011111000011001000010101010001111101101010011100000000110000001011100; 
out3768 = 128'b01000000011100110100100001011101110100001011110110101011100110010001110110000001100110101100111001111101010110000001011011000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3768[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3768, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000011000011010001011101010110100011101111000100000100011000001110110100000100010101101101010101111101000101011110100010101; 
out3769 = 128'b01111111101011011101000000101010100101100000101100001000110001100100011100011111011001101011111101110000010011000011101001011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3769[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3769, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000100010011111100101101101000110111011000110111101011010100000101110000101001111011110101001000101001001101010100000101001; 
out3770 = 128'b01110100110011001100010010111011011111011000000011000111111101111110000010111101110001110111010001110001001110101001101111001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3770[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3770, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010100101100011100110101001010011010111100000001111101100011111101010101010110010110100001010100101000100001011100011111000; 
out3771 = 128'b00100111001110011111110011111000011110011101000100101111000001011010111001100100100010010000000101111011100011101111011000110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3771[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3771, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100001110110000001100101110110010101011001010100001100111111110010010101001010111110001110011100101101100011111011110100001; 
out3772 = 128'b11011110110101110010011000110101010000001010000101000011111110010101110000110111010101011010111011111100101110001111011001011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3772[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3772, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000011111111101010100000111000111110011110001000110110100010011001001100101000000111110001011001100011100011100110001000001; 
out3773 = 128'b00001101011101101000010001101011101010011011010010001100111111111000101110001111110001111101010110000010011011011101100111001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3773[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3773, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011101010100101010111001010010000011110010110001111111101110000100001000111110110111010101011000110110100100111001100011000; 
out3774 = 128'b00001101101011111010111011010101111101011101101001110011101011100000110101000111001111011111011001111010100110000000100111101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3774[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3774, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110010100001010000101010011010001001111100010011001101010001110001101110101001011000111100000111111110100100001011110101110; 
out3775 = 128'b11101011001011101101110110010001011101111000101110001010000100001010111001100011010010000100000011101101001110011000011110010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3775[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3775, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101111010001010110101100100100101100100000100111111110000110000111001101101000001010011100000100001011011111100100111001100; 
out3776 = 128'b01011001001011110010001111101100110011111011100010001011100000000011001110101100011000010100111010100100111000110110101011110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3776[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3776, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110010011100010010111111111010110000011000001001000110101111010100101010000111011111111011100000001011001001010110011100111100; 
out3777 = 128'b01111001010010101010001011101101001010111100001011000100001100110101101010000000010100001001111111101011011010001011100011110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3777[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3777, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110000010011101001011101010010100011010110011111000111100111001111111000000101101100010000010010001101111110101111111101111; 
out3778 = 128'b11011110000011000001010001100110110101111111001011101001000110001111101010101011001100100000000010110100011001110111100011111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3778[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3778, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110101100011001110000010010110001111110110100011011000001100111101000000101000010110111100111100110111000000011001001010000; 
out3779 = 128'b00101100110110100010010011101001100011100101010011111001100011000110111011100001011000001100011011100100100001100100101111100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3779[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3779, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000100010101100110001000110100001101011001111001111110110110010101000101010011011010101000010111011100110011010101100001100; 
out3780 = 128'b00111110011110001101010101001110010111000101110010011011110001001100100001001001111111111001011010100010110111001110010101110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3780[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3780, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101100010010001111011101011001111100100101000011101111100000100000011110101101000011110010000001011001011011100011000010011001; 
out3781 = 128'b00100101001000001111011101011111111010001110010111110000001001000000011001011101010001111101010000001101100110010010001011001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3781[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3781, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111011110001111011001010001010100011110011011110100101010110010110101101011100010110001101001100111000000100110110011111110; 
out3782 = 128'b00110010100111101010000100100110111001001010001010100110000111001011101101000010001000101010111010010111100111000110100011110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3782[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3782, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110001001111100001000110100010100011001010111101101110010001110110111001101010110111111111010110010111111011010110010000001; 
out3783 = 128'b10010100111001011111111001011010010010100011011011110111010001011101110011111111010101101000111111010101000101000011010010100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3783[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3783, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000000011111101101011110100111001000100001011010100001110100010000000011110010001011000110000010100001101111100111110101111; 
out3784 = 128'b10101001011110111101101100111010001011111100001101110101011100110000000111010110010101001000010010010110100100110010010101001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3784[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3784, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001101110011111111101111100111010001111110100001000000100100010111010110101100100000000000101001100000111011111010001110110; 
out3785 = 128'b10101000111010010001001100011010010000100010001111111011110101001001010111101011011000111111011010011100111010010111111111111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3785[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3785, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101101001100001001101100011111111011011001000001101100000000101111110010000000011111011010000000110101101111111011111000001; 
out3786 = 128'b00110010100111011011000110010001011110000000011010010110000011101000011000111111010101000100101001011011011000010111000001110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3786[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3786, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000000000010000011100101101110110000001000001010010110110010111010011101001110011110000011110100100100111011011010011010011; 
out3787 = 128'b01011011111110000111001101000101110010010100110111101110000110110000000011111011111011010000111110101111111100000001101110011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3787[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3787, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110000010011101101000000110001010110001100110010110100110010101000011000000101000011010100110101001101001111011010010101011011; 
out3788 = 128'b01110111011101101001010010101101100101110100110010111110100111001111010101101011011111101101111111100111010101011100011000111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3788[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3788, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111101000101101101011101111101111101110101111010111111010001000001010000001100001101100011100111000111110011111101110111101; 
out3789 = 128'b10110000001010110101011100110001000001100001110101111011111011001011110101110101001111010110011010011011001110011110000110011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3789[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3789, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011101011101000110001000010001111001110100000000100101010101111111100010010101101010111001011101111100000110111010010101111; 
out3790 = 128'b01001101001011011010110010100001001101100101011001111011001101011100101000110101100011111001010110101100010011101111100000101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3790[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3790, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111110000101101000010001100101111010111011000001111010100011001111111101011001010111101101001100011111101111101010101110101; 
out3791 = 128'b10000010000110100110011101111000111111101011011100101000101011110100010000001111011010101001001100010010100110000001101001001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3791[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3791, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110011010001110011000111101101010100001000111111101001110110100010100011101010101110010011010010101001111010010000110010111; 
out3792 = 128'b01001011001000011110101111011110011010100010011001001111010010110101010111011010010001010111111101110100101110010001110110100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3792[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3792, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111011110110100101100011000111100111111101010101111100000001110010100010101101111000101010100011011111101111010101101010010; 
out3793 = 128'b00101000000011110110111100001011101111000110000100011001110011100110001001000100111011111000111010011011011101001100000011111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3793[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3793, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001110101101011110111000110000011000101001111100111000100010001101110000010001100010100100001100011010111111000101010001000; 
out3794 = 128'b00010011000110101111111001001110101000000111111011010100000111110010011011001011011011010101110100011011010001110001000111111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3794[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3794, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011110001000010110111001111100010010001100111110011000000100001100011111011011111101000000001100010100111001101101100010101; 
out3795 = 128'b11011101010111000100001100110101100011011011100011110111010100110011001010010000011100110101011101010010011100001011100111001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3795[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3795, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001100011010110110010010000100010101001101011111000011110100010101111110110100011100001111110010001111100010010011000011001; 
out3796 = 128'b00110000101111111111001101101001111111001001001001111011111100111001000001001111111000000100100110010100111010000011001100001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3796[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3796, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100011001101000100100111111000110001000010000010100010011011100100001011000101001101100010101001111100101110101000001101101; 
out3797 = 128'b11011100000010110010111011000100101100100101000000001010011001000001011100010111110011011000001010010000010011000010011011100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3797[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3797, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101111101100000111101000001101000110110100111100011000101001110011110110110010001110100010011100100110001010011100110010010; 
out3798 = 128'b10111100000001111101000000101101111111011001000000100111101011100100101010100000100111100101101010101100101001011010010110000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3798[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3798, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101000000001001011000010101010101101101001001101010000010100001110100111101111001110000011001001110101110110111000011101110; 
out3799 = 128'b11100010000101111101010001111110100000001011101010110011111110010011000010111011000100011100010110010011100010001101010010011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3799[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3799, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000100000100001100000101111101011010101001110011000010100000100011110010010000100100100001111011000011110001000101010001011; 
out3800 = 128'b01100100011011101111110111111110011101010001100000100011111110101000000111000010110101101100000100010110100011111000010010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3800[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3800, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110000110101011010010011101111010010110110111000011110111010011111101100000011011000010001100011000100100101101001001101101; 
out3801 = 128'b01110101101010111011110110100110010101100110110010101111101011111101110100100110010110111011100011000001111011111000010010011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3801[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3801, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010111111000011100011010101000111111110101100001011111101001111011111011110101001011100000011100100100110111110101010111100; 
out3802 = 128'b10100100011001000011111111011111100001101101111101110010100111111111111001100111101011110101101100100100000101000110101100110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3802[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3802, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101000001100110100111100100101100000000101111110001010110101111010111100010001001110100100110011010001101010000110000100010; 
out3803 = 128'b01011001011110010100111010101001001000101010000000010101101000001001000101001001110011101110110111001111001011010000011101101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3803[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3803, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011111100110001010101011011100100111001100011100001001110100010111101011000111101110101010001111010011000011110000001001001; 
out3804 = 128'b10000000111010100100110111101001001110110000101100101111000110101000101010011100010101101111011100100011110010011011100111101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3804[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3804, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100110110011111001010011101000001011100001010111000100001001010010100011111001110010110110000001010010001001010011001110110; 
out3805 = 128'b11111001000010001010000110000100001100000100011011010011101110010101101100100011110111011111111001010001100011110000111100011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3805[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3805, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001111010010010111100110101101001110010100111010101001100110010100010001100001111011110010000111010011101000011010001111001; 
out3806 = 128'b10101111100010011000100000100100001101101000111011011110001010011100000100100101110110011001110111001010111100101100110111011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3806[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3806, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001011110000011111001011101001000101010010111000011000001100001110101001101010110000101111111000000000010011011100001110101; 
out3807 = 128'b01101110101110111111110000001110010001001010111001000110101011111100011000010000011001010010101100101111111010010000101111010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3807[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3807, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100001000100011011100101010110110000000000011000111011011100001111011110001100111101111110101110010111010101110101100100011; 
out3808 = 128'b10011001010010100101001000011000100000111010000110100011100010000010010110101111111110100111000001100001101100101110010100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3808[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3808, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010100010101011010010000110110100111010010010010110100101001000101111110001111100100011100100111110001001110011010000100110; 
out3809 = 128'b10111100011001000000101110101110110110011101110011001100010001011101010100100101111111000100100011000100001011011110000010110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3809[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3809, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111001111000101011000110110100101000011001110000001111101010111001111100110110010010011010001111100101110100100110111111100; 
out3810 = 128'b11110100100011010101011001100001100100111011100111000111110010100110101010010101100010011100000110001111111110110011101101001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3810[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3810, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100011001001001100110001000000000010000001111100111000101010110110100111001100111101000001100101101111010111111101100111101; 
out3811 = 128'b01000001101000110111010001111010010101010011110101101010100011100100001010010111010110111011100110000110101101001111100001110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3811[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3811, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110010000001111001100101001010010010111101100010010110101010100011111011111100011101010010100000011011000001110000101010001; 
out3812 = 128'b11001110000111011111000001011010001000010010110110010001010001010101100101110111100100010010010010110010101100101100111011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3812[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3812, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100111100011000110111001000011010000111011110011011000101110110010111100111110101101101010010111101101101110000111100100010; 
out3813 = 128'b11111100011110101110011001011101011111001011110110000001111001110111101000100001001111011010000011001011010111010100111010110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3813[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3813, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000000001101010001110101100101100010001000010110111011101111100100001001000100111110000111010111101100001100100110101011001; 
out3814 = 128'b01111100111011100110110010010100001100011100110000101010110010011110011000100011110101110011111100000011101010000101010010101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3814[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3814, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000100100110000110000000110000001111001000001110110101100001110010110011101001011111001110110110100001010001100100100001001; 
out3815 = 128'b00010111110100101100110110101110001011001011000001000110000011101010110000000111011110010001001101110111000110111110010111100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3815[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3815, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100111001100010110011101010011001110100011001010011011110010100010110011111110011100110000101101100010010110001000110001011100; 
out3816 = 128'b00001100011011100110101101100101000111011000001010110101010000001000100010101101101001111100010100010101100100000000101111001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3816[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3816, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100000100000101001111001100010100010010010101101000100011110011000001110000111110000111101011100011110110000111001001101010; 
out3817 = 128'b10000111001011101111100110100110000101101110000101000111000001110100010110010111100011001001110110001001000110001010011011100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3817[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3817, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011100010000100001000101111001010001010000000010010011111010001100000110011111010100100110000000101100010101110001000011110000; 
out3818 = 128'b01111110001000110010011111010110110011110010110010001001111111001010010100100110110001100011011101101110111101011010111111011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3818[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3818, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101100101010011010001000110111001110000000110111010110011100001111010110011110101101011100010110101010111001000000010010111110; 
out3819 = 128'b11101000110101101101100101000000100101111010000100111101100001011011010000101111101001010000110101011001001000000100101110011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3819[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3819, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111110110011110110101101010000001001001101110000101001100001100101100000100011011111001011001101010110100101110111010100011; 
out3820 = 128'b11100110100110110010100011001101010011100110110100110010001000100110111100010011010111010111101101000100010111011101010000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3820[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3820, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110001101010011000010101101011001101100100100110010100110100001111100111101101100011100011001110010001010010000010101110101; 
out3821 = 128'b00010011010110110110000000001010101101100110100111001110101001100111100111100011110000101001001110100100100101100110100110000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3821[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3821, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010010110111110011010011101011100110110000000100000010011111011100011001011111011100011110010111111110110001010010010010101; 
out3822 = 128'b11011101010111110110111111111111000011100010011101111101110001111001111000001010101011001000011110100111110000000011001010111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3822[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3822, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001110110001011110101111001011110000111010011000111100001100001001101110001000001101100110001001100010010011001100010011110; 
out3823 = 128'b10001001101101101010001101010010100111001001011110110111101001111101100000110100110001101101110110000001001011101001000101010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3823[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3823, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110000101111010110011111110011111011111111011101010110010110000011110100111111010011111101010011111111011100110101001100001; 
out3824 = 128'b01000101101101101101010001101000000101100110110101000101110011010110011111101101001001010000101010000111000100111111000010000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3824[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3824, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111110000001101010111010001111101011111011101110011011101100001001100111000111000100010000100111111010010011001100110101010; 
out3825 = 128'b01010101110100010110101000011110101010110000111100010010000101101111000011110110111100010000000001000111000000111000110011010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3825[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3825, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000010111101001010011010011100000011011000101011010110101001000011100000110101110010101011011001100011000001110011101111101; 
out3826 = 128'b11111001110000100000010011001100001101101000111101000101100010100000010000101110000001000101100000011010101010111110010010111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3826[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3826, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111100100010101001001001111110000100000110000100001011010000011001011010111110000100110011010010100011100000000101101000110101; 
out3827 = 128'b00000100101101111010110000110000010111110111010100101010101011000001111111010111011100100100100000000111000010100000100000101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3827[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3827, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110011101111110001001010001101100111110100111000111110000111111001100111111001100100010011011100100110001100000110010111001; 
out3828 = 128'b01001101000011001110101011010010101001001101101000001001011011110101100001101110100100111110011011001010010111011101111111000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3828[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3828, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101100001111011001000100101010001111101110111000100110011010111100110001001001101110101011101100111010000011110100000101001; 
out3829 = 128'b11110100001100011010000001010011100110010001110001100100011111110100101110010001011101001011110010010000101001111101010010000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3829[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3829, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001100011100000011100010000110010001010011011101111011010101111101101000011100100010101010000110110100110101100111111110100; 
out3830 = 128'b10001010010101111010001101110111001010011100100000100001100011111111110000011110110001000011111100100100110001011110101110001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3830[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3830, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101100101001000000101000111000110010000101001110000001010111010001110101110000110110011100010001100111011111100110001000001; 
out3831 = 128'b11010111111111101110000001100010101010101100000010010011001100001011010000111101011001000110000011010001011100110000100100010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3831[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3831, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100110010010001010110111011010010000100010111010111000101111110001000000110101101001001001011110011011111111011101011000000; 
out3832 = 128'b00001000000110010100011010000000110010101001110001011100000011000111110011111011100010101101111100101100011001111101011000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3832[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3832, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101001011111010000000000110101000110000100010101011001101110110010011111011111101001111101001001011101101111010001000001110; 
out3833 = 128'b11010100111010101000110101101111001110010100101000101110100100011101001011011110101110001101111010011110100110101011110101101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3833[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3833, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000011001100111000001001101010111110001100101010010000110010000001010010111010001011011011001111111100000101101111011011110; 
out3834 = 128'b11111111011001110010011000110011000000011010101011101101111010000100100111110101001000000011000001000011010111001100011000100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3834[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3834, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011001111000100000010011000010100000001011111111100100000011100111100110001100100101110001111100110101101110100100010000100; 
out3835 = 128'b00100010010000001110100011010100110111111001011111000100101011011110001101010101001100011100011010000010111000110111110101011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3835[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3835, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110000101111000101001011110000100010110010110010000001011101011010000111001010011110000011011000010110011011101111011110011; 
out3836 = 128'b10110100001110100001011101111110000000001001010000000101111000110100001100101000001110101000001001111000011011011000111100101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3836[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3836, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111101010010100110110000000010001111000100101101101111100111011111001010110001000111101010010011110011110111110011011110000; 
out3837 = 128'b00011100100011000000001011111101001000110000001000111010011000011100110101010111110010000000010001011110001010110100010101101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3837[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3837, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101001111010010000011000110010000111000000110111111001111110100111101010100000011100100111000101011110101100001001100101010; 
out3838 = 128'b01111001000110111001011011010100001110001011101110110101111011101001101001100100110101110010001101011101001101101011011001110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3838[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3838, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001111100101101111010101011010010100110101011111101110111110000110100110101011101110110110000010101100000101111101011100101; 
out3839 = 128'b00010111110001100101001011000010110110101110011110001100010111010000010111010001110010001100000101110110101011100010110110010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3839[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3839, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001011010110001100010000110110000000101111111110110001011110000010010011010010100001111101000001110111110100110100101110101111; 
out3840 = 128'b00000001100110111001111000110010111101101111100001010000101111000101001000010001001100110011011011100001100110001000011000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3840[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3840, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011111010001001000010101010101100111011101001001100101101100110010100000010001110110010111111100101110011100000011010110111; 
out3841 = 128'b00000101101010110001110011000111010110001010010010101111111110001010111011001110101000010010001001000111011010000000010110000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3841[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3841, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101110111101001100101101101010000011000010100101111100100110010001101000100011111011110001100001001010011010000010010001011; 
out3842 = 128'b00011000001010101110011000000111101000111110110011101000110010001100011000000110111001101001110101101111011110101101010100010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3842[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3842, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100100011011101010101101000111111101100111100011000111001011000101100100101010101100101011101010000011100001000010101010000; 
out3843 = 128'b01001011011010011001011101100110010010011110010100010101110100001101000010111010010010100111111111001101110101111100110100100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3843[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3843, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111000010101100111110100111111010001001100000000010101011110101101111001111101011111001100110101011111001010110101001110000111; 
out3844 = 128'b00011100101101101010010011100001011101101000000001011010010000000000001011001100100001011111001000011001111110110011101100000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3844[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3844, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101100010001010010110010101001011101000111100110011111111100111010111111011110001101101110010000101000110101010001001000001; 
out3845 = 128'b10000000001100100111000111010101001111011011011111011110101000010001101001011111100101101101101000110111101010101011000100110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3845[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3845, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010100010100101010010001111011111100001111110100010011001101101111110000111111101110110100000101001000011000010101101110000; 
out3846 = 128'b11001010001010011100111010010111011001111001101010110001100110100111101011010011011110111100001111110101101101110011001101010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3846[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3846, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100100101000011101111011100001110101011110100011011011011001100101010111100011111010001101000011110100000110000101111010010; 
out3847 = 128'b10111111000100010110011010101001100001001111001011101010110001010000011011110011111100111111000100001111100110101110110100011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3847[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3847, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011101111001010101011111000101010101100001011100101101010100001110001111010111000001100111111011111111101111001110100101111; 
out3848 = 128'b01011111001110101100011111100111111101110000101111010000111001101110000011100100000100100110100110000010001110100101001110110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3848[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3848, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110010111010110101001001011011100000110110000101001101111010110010101110100101011111100010111101001101100001001101010001101; 
out3849 = 128'b10110011101100010101010000101010001010100001111000000101111010111101010010111011111011101010001110101101010011000001000001110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3849[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3849, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111100000000011110111001111100000000001011110111000000100100100010110111110010110010011011110101011110100001111011010111001; 
out3850 = 128'b11110111001010011110010000011000101110111100100110110101110001111111111100110010100110101111011110110111100010111000011110101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3850[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3850, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110101010011101111000000101000000111111010001000001011010101100111100010100100000111101101111100100001000111110001110110010; 
out3851 = 128'b10111101111111110010100001111111101101101000010110111101101000111110110011010100110001000111111100011101100001000100011000100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3851[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3851, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011010000110001110000010010100100100111100111001111110100100010001101001100011101111000000110001011011100000000101101110001; 
out3852 = 128'b00001000101101011111010110011010111001011000111100011011010001110101110101100110110010110001100111000110000110101100101100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3852[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3852, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101010011001010001110100011111101101000000000101111101110001000011011100011000111000111010100111010100101000010110001111100; 
out3853 = 128'b11100000011010001110111001100000001000010000000010101101000010001000111101111111010011011000010000011000110111101000011110101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3853[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3853, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100111011101101001110011101001110101101110110001011101110101011001110011001111110100011100010100000100101010101001110001100; 
out3854 = 128'b10011110011110110110010101111000100101101011101001111100100101010110001111100001101010101010000110001111001101100110100011101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3854[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3854, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100010111110011111111010010100101010111001101111100101111101110000010010101101100110101001000001011110111001011100110010100; 
out3855 = 128'b10011111111010001011101101111100101111101100010111010111101001001010111001101001101100010000010011001000011001001011100011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3855[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3855, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011001111011100110110110111111101010000101100111101111101000000010110010001101010011000101110011000100000000000011100100001; 
out3856 = 128'b11000000011100110001100101011011110001110101110001000010010101010101110011011100001101111000101100011101101110011011000110110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3856[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3856, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110001100111111001010000111101011011011100000111101100111001100000101101001110101100100101110111111110000111110100000000100111; 
out3857 = 128'b01101110100010101010001010101111111011111011001001100000010111001010110110000110111011101010101111010000001101001000010100101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3857[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3857, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110100100110111010101100010000011001011000110110111011000110101001000010011011100000111010110000010000101011011010110011101101; 
out3858 = 128'b11010101100111101111111010000100111101010010101110000101111101001011000011110110000000100011000110111011101000101110100110010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3858[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3858, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010000001111001001100011010100010111100110101001000011000111000111011110001001110100011101111000110001001110101000001010110100; 
out3859 = 128'b10100011011011000000010001101110010101010111010110000110001111100011011100011110110011101100100111001110100000111000010001100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3859[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3859, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100111010101111100000101111100011110101010010111110001001101011110100010010000110100011110100111011011111110111000111010010; 
out3860 = 128'b11011010001101100000000110011001100010010001101000101111100001011101010000110110010000101001000000111000011000100011110010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3860[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3860, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000110010011001111001100101001001000001111100011010111011101100010100010100111110110000100101111100010110011001101110000010; 
out3861 = 128'b11100001010000100010101010000100100000000110011111000100011100101101010110011011101100111011100100010111000011011101011111111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3861[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3861, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110101001011101110110110001001100100001011100011011110100100001001001111111010010000110101100001011011100001010101001111000; 
out3862 = 128'b00001100101110100000110110111000010101011011011011011010110110110111000100011100011011010011000000100010101010111101100011111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3862[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3862, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100100101000011110010100000001010001000001001100111000001010100101010001010100000010010100011001111011001000001011011101111; 
out3863 = 128'b01101000111101001110001111000101001101100100110111011110011100111011011101110101011101001110011101110001011101110110101011101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3863[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3863, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100100110010011110000001011010001011010011001010000101100010101011000001111110111000101101010110011100011111010101101110000; 
out3864 = 128'b00011010001000100011101101010110001001001001100111111010101101101011001100010111011100010111000011001101110111110100110110001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3864[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3864, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101000010111011011101101100011001111010101000111010111011100010101111011001101111100000011101011010011111010011110010110110010; 
out3865 = 128'b11111101110110111101100110010001001001100011100101000011100111001100001001010100100000101001010010001000101010010010110001000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3865[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3865, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111000100001010110010110110001001100000011101000100011100111001001101110010011110111001100000000110110011011001010001111000; 
out3866 = 128'b11101001010001011011000110011100111011001010110000011001110101111010101011111001000000011010101000110111110101110011000010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3866[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3866, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011010011000101011011110010010111011100011111101111011010100111101100101011111000110000010010000100111010011000000100011010; 
out3867 = 128'b10001000011110001110010100111101001011101011011000110001100101111001100101110011011100010100111110010000001001011011101010001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3867[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3867, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000000110000001011001100110000110101001110101111011000011100110010101111101101001000001110110111101001110011000011010011111; 
out3868 = 128'b01010011010110000100101001100111011000001111000100010010010111011101001101111110111001001010111100010101001001000001000111101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3868[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3868, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000011101000011000101011111000010000010110000111111000101110010010100000110111000001111111011110001100100011011011100100000; 
out3869 = 128'b01101001111100100100000100011011000111000001011111100010001110110010001010100001001011101001011000110001110011110110100010011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3869[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3869, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011000111101110001100110001110001100001100111000100100110101110111100011001110101111001010110000100110111011010010001001101; 
out3870 = 128'b00010001010011011111001100000000111101000000100001100110000010000110110100111001000010100101010100000101010110001010011010101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3870[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3870, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000111101011010011100101010110001101010000110010011101111001101010100011110010101100101000001010110000000110110010000100100; 
out3871 = 128'b00101000000110110010101000001011000010110111110010010001101101011000010010100110111000001000000001000011101000011010000011110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3871[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3871, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000000110110111101101110001011001010011001010110000011001110010100010100010011010001000101001011110111111100100100101110111001; 
out3872 = 128'b10001001111000010100001111000010011000101000110000110100110110110110000101001001000110110101111110111100100000010111110001000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3872[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3872, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000100001101000100111101110101100011011101101000001000100110110111000111001110000001110100100001011100001111101100100011101; 
out3873 = 128'b10011011011011000011011011101010100001010100100111001100001101110011010111100000100111011010101111100000001011110110001010011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3873[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3873, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111111000110100111101010100000111001110111101000100100000101110011011001101001100100000111110111011110011010010101000111001; 
out3874 = 128'b10001010101111010111000001110100110010000100110101111111110010001101000010111010111100110011110010110100011010101111101101111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3874[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3874, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010011001000110110011111111111001101010110110100011110111000000101010111000100110001011111100110100000001100101010100111011100; 
out3875 = 128'b11111001111111010110111110110001000011000010111001111100010011011101011100011011010001001111010010101001110100100110101001100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3875[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3875, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101001001000011011110100011000001011001101011111110101011101000101011011001000101100100000110000100001010010100111101101110; 
out3876 = 128'b00001000111100001101100110010100001101100110001001011111010101101001000100000001011100011010100100000000011110100111100011010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3876[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3876, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110111110000000111111111010101111101000100110001101100111111111110001110111000111100000010011110001110010000010001000111000; 
out3877 = 128'b00000101100011010110010000110011001011001100100001101111101010110010010110111000000001100000011000110011101010011100100110010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3877[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3877, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011000010000000011111111110110111111100110001010111010100110100111100010011110101110001100001011111101011011110000101010010110; 
out3878 = 128'b00000010001101100111101110000001101110110100111000111111011001010100110010100110110110010011111111011111111001000111001011010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3878[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3878, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100001011011110110000010011100010110101111010111111010101001100101111010101100110110100100011010111000011101010111100110001; 
out3879 = 128'b10111101110110111010110000001011111110100110100100100011001100011011001100001100001000111000111111110111110101001111101010000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3879[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3879, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100100111101010110101110011110110111100000110111011001111100110100011011001010000110000100001100011011000001011100011100110; 
out3880 = 128'b10000001001101011010100111100001000101101100010000111000101111110001110011001101000110110010010000110110100111110000011010111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3880[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3880, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011001011000000101100101101000011101111010110111100001000011110101011000101111000011111010101100101010001000001100111111111; 
out3881 = 128'b10110001000000100001111101101110101111000110010101000110000101101011101011111101000011111010011001110101010101110001111010101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3881[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3881, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101111000111101100111101100010011011010100100000100011010100000011111101000010101100010000111010111011110101001011100101000; 
out3882 = 128'b01000100101100110000101111000010100000001110011110111000100001111101101011010111010011000110011100111111001100000001101100011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3882[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3882, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010011110101001111001100010101111001011001110000110100001000010100000000111111101001111000110111001001001001001111010010010; 
out3883 = 128'b01101111110110011001011011110110101110011011011010101010011011101101011011111000000001101100110110010110101101100010101101111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3883[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3883, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111000010000011100111000101100101101010001010000110001111001110101011000110011011000111010110010010001000010000100011110001; 
out3884 = 128'b11100001001010111000111010011110000010110001000110011100101111101011100010111000000011010111100000100010110111001111111011111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3884[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3884, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101101001010010010001000011000111011010111111100010110011111001000100111000000110110011000010011000110011010110111000111101111; 
out3885 = 128'b11000010011100111101000110110110101101000110110100101001101010100010100000111010100010101001011101000110111110110011000101010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3885[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3885, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100000011111100001000001011101101011110010010001011100011001011111101100000000001110110011000100001101001110100001010010000; 
out3886 = 128'b01100001110001011011111100100100011111110001101110111100000101000111000000110111010101011000000110100111011111010000100100011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3886[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3886, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011011010001010100001001000011001111111101001110001010100000001001100100110000011100111101111000010101001010011101001100011; 
out3887 = 128'b11101001110111011111100101000011111010001011000110001110010100011111101111010111101101010111001000010100100100001000010101001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3887[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3887, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101000100010111110001010001101011110001110001001100111010111011100100101011011010010110011001001100100001111111111001101000; 
out3888 = 128'b10101110000111010010111001011110111101000110000011111000101000101010101010101111111111010001111010010001111100001000010100111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3888[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3888, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100100101110111010010001110110110001101001100001101001100010010100101001001100100100000111010010101000111011101001011110111; 
out3889 = 128'b10110111000100110100011110001100001000010110101100111000110100000010001100010111001001001011010010111011010100001110110010111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3889[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3889, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101111100000111111011000010111110101010010100001100110011000010001001110011000101011110111010110101110110011010000011010101; 
out3890 = 128'b00011001101011001111101111011100001011000111010101100011000010101011101010100011100010100101100110011101010001001100100000101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3890[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3890, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010000110111001101110101011011110010111101000011110101101101001110110011000100110101110110101110111000010110110111010001000; 
out3891 = 128'b10111111001101111010011100110101101111100101100010110000110000100110100001111010101000101010001001111111100110010101101001010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3891[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3891, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000011000000101101111001000101110101000010100011110010100111110100110001111010001110001101110011011000010110010101000111000101; 
out3892 = 128'b10101010010110100101001100100111000110100000000000111100000100101110001110110011000101101101100011100110010100100101011110011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3892[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3892, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001011111000101010101010110101111001110110110100010000100111110110001011010110001010100010011001010110010011111001111011101; 
out3893 = 128'b01110101000111110111101101111110100111111001100101110010111000110110010000011001000000100011110100100011110001000001111110111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3893[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3893, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100011101111010100001110101001010000011100111111100110100100110111111101010111010000110000001100101100110010001111001101000101; 
out3894 = 128'b10100101111110110001011001100010101010001100101111011101101000111101100101101011101110110100110101101010001110000100101011100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3894[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3894, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000000010000111011100101001010110110100001110100111001110111010011010100011111111111001111110010110101101000101011001011000; 
out3895 = 128'b11110011010011101100010111011001001100100000110001001110101000001001011001110111010001101011111001111101101000110010001001001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3895[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3895, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000111110011111111000000100010010001101001110000110001111010000110001001001000001010100111011000000010000110110001011010111100; 
out3896 = 128'b10011100000011001100110000011001000000111110010011001011101010001011000101101111110101011111011110011001100010000010001111100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3896[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3896, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001110001111110011111001011111110010011000101111101011110000010001110111011010100111001101110100111111001101010001101110110011; 
out3897 = 128'b01011000010111111111010101101010110001010000000100000011101000000111110101111111011010000111000111001011110010001001001000110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3897[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3897, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000001001110111011011101011101011011010010000010100100001100101111100111111111110011000101010000011111011011111111110110000; 
out3898 = 128'b11110100000101010011011110100101001010100111001111110100010001010001110101000011010101000000100100100001010101001111011100001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3898[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3898, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111000100001000010111101001100110111100010011011001101101000010001010100001101011011010011111110011010100101001111001101110; 
out3899 = 128'b10001111010101010010110101111000010011101111110001100011011001100001011010101100111110000001001011000100111100110000000111110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3899[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3899, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011011101101000001110100010110001110011000100001001110100111101100001101010100100011101100101101000001111110000000110100111; 
out3900 = 128'b01110010100011010000110110001011110011010111100000101100001110011000111100110110101110010000011011100110110100100111110101011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3900[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3900, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101110101011111011111100000110100010111100111110111100111011000110111110000111000111001110111101010110110011110001100110011; 
out3901 = 128'b01111011101000011011110001011101000111100000110011011110111000000111101000001101111011111001101010111101010101100111110110010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3901[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3901, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101110001110010011001010111110010111100000000010000100010010001001000001001101101100001100111000111011101100100001001011101; 
out3902 = 128'b00010010101110011010110000010101010001011001011010100111010010100100001111101110010010000101111001110000010101100010000100110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3902[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3902, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001011111000100011101110100011001110011010000100000100110011001000010001011101000101010110001101001100101111000110000010000; 
out3903 = 128'b10100101001111101001111010100001111001111111011001000101010011011110111000000110000011110000110001001010011111101011110111000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3903[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3903, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100100010010110010010101101101001100101111110010000111100010111000101001011010011001011011111110100100001000011111010011011111; 
out3904 = 128'b11011010100000101110110010011011001101100000111111100000110011100110111110100001000010110111111111010111101000111111010111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3904[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3904, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010101101100111011101101001101111000011100101010110000011011001100100100101111100100000000101100100110010010000000100010100; 
out3905 = 128'b10011010010100000100010100111001101001100101101100010000110001000011100001100111100111101111111011000110001000100101000101110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3905[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3905, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000011000101010111011110111010101111100011010001011110011010111000101100110001001000001111010101101100100001111111111111010; 
out3906 = 128'b01010111000111111000011111011001111110100111011011010110111110011010010000111110101100000100110000100111011111111000110111011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3906[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3906, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000011111000100111100000101110100100000000001100011011010000100001001011011110001010111010100011001000010100110011001010011; 
out3907 = 128'b00101001100011101010101110000111101100100100000100101100011000111010011110010110000010101011001001110010101001110111110001111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3907[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3907, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100101110111110101101101111100101011010110111001001101110110110000110001010111111101110010100100000111010110001111010101100; 
out3908 = 128'b10010100010001101001000101100010111010101100000011110010000010100001110011101100001111000000111001110010010000000000101110001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3908[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3908, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100000001110110001010001101001100111001001110101011000111101001011011110011111000100110011110101001000100111001100011110011; 
out3909 = 128'b11100010010111110101100100100000010100101011110110001100110110100011011010111001011100100100011001001010000110110110010111100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3909[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3909, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011010000100001000010100101011100010001001111110110110111011011010000011001011110011011001000100000110111100111111010110000; 
out3910 = 128'b00101101001011110001011111100010101100011110101110011101100000111100001011011101000000110100110010010011110011011011111100100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3910[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3910, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010011001010010110100010111001011110010110110000100000000110001100110100100010111000111100111101011010100001110111001010110011; 
out3911 = 128'b00010100000001111110001101101100101000101101001001010010111110101001100001110000010100111101010011110100110010001010000101100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3911[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3911, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100100111110111011001001011110100001010000001101101000000100101100111001000001011111011100010010011111100110111110011011110101; 
out3912 = 128'b10000100111000100000010111001100011001110110101100001101111110100011101111110001100101001101100110100110001011111101001110111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3912[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3912, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000001000011001000010000001100001000000011111011011100110100011000011000100111100011010110101010110010100110001011000000101; 
out3913 = 128'b10011101010110111010010100010101111101010001001000110100101111111011001011010011010100100111010111010110001111000101100011010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3913[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3913, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100000011000010011010111010000110101001001010110010110011100110011000000011010101110000101001100101010110000011011001010110010; 
out3914 = 128'b01000101000101000001101011100110101101110111001000100000001001110010111000000111000100000101111000111101101010101001010001011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3914[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3914, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100010011101110000011110000001011101001100111101101110110011001110001010101000010100000011111010011100110011100001110110100101; 
out3915 = 128'b10010001011001000011001100100001100001000101110011000001111111001101110011011101100101111101101011111001101100001011011011001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3915[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3915, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101000001100001101101000101110110110000111111101001010101010011011010000111110011010010011100001000111111110111110100010011; 
out3916 = 128'b10101000000101111001110011101110001101001000101111101111110000001010000001001100001111110111110001111110111110001101011000000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3916[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3916, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100101111100101010011000000000110011110100011010001001111111010010110100110010111010100100010010010111100110010001000010111110; 
out3917 = 128'b01101001011100110001001111001000111101001011111000010111011010100011101001000111111101111101000010101001001000010100111110000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3917[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3917, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000111011110110010001000001001010011000111010100011000011001001000111000001110011000001001001001100001101111010111000001110000; 
out3918 = 128'b00001111001000100001100011010011000101000010000111101000100010010000000010000110111001110000011010111100010111101000001001101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3918[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3918, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101101000010000100010100101000001101100010100100111000010100011101010010011010001011101000100001001101110010011100011010011; 
out3919 = 128'b01010001110010101001100001011110110111001101100000101100001110000100101000100110100000101101100011101100000011010011010001110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3919[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3919, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011110111100101101001011001001010111110000100011010111000001000010001001000111100100111100010011001001011111110011010000101; 
out3920 = 128'b00000011110000010010101101111011000011011110110001100000010000101111000100001110101110101110011001111010010010101000001011100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3920[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3920, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110100010111100111010010100000000111101010111001000000111101101000010111000001111101111001000101101011100101100010111011100; 
out3921 = 128'b11011010010111011010100101111010100011101011100001011011101100001110100111011010110111000011111101110101101001100001010010111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3921[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3921, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011111010101100100110111110001000010100110001001010010110110101011001000001110001101011001101101100001000011100101001011110; 
out3922 = 128'b00111100111111000110101101010110000100001111110001011011011111110111100100001010111110110101111001011011111000111110011010001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3922[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3922, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011000111110101110110111100000000100010001101111011000010101001000100001011110100101110010010101010100111001011011101100000011; 
out3923 = 128'b00111111011001101011111011100101000010010111110010011111110100110101000101011000010111011101011111000000001001000101101100010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3923[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3923, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010001011100000000010001010011111101010100011001100011000100110111100110100001010000001110010100101101000101000110101111000; 
out3924 = 128'b01000101000011001001110110001110110000011010100011000011100101011101000100101001111100111100101101100001101100001001011000101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3924[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3924, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000001011000000010000110100110111101001011000100111111010000001111001111000110111111110011111001100111111101001101101001000; 
out3925 = 128'b00100000110101010110011101111100010110110000111001100110001011100011111101011100110000011101001110111100000011100101111001000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3925[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3925, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011110111110011000110110111001010011100111001011100011010101100100100001000001011101000010000100000110101111101001000011110001; 
out3926 = 128'b00011001111010000000111101000100000111011001010010110001100010111001110111100011111001101010101010011011110000100010100000011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3926[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3926, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101001001011100001000110000001010111101100010111100010101011010110111000110111000000010110111011001000001111001101110110100; 
out3927 = 128'b10001011110011000110000111000010111001010001000110101001001101010100100001111010011001111110101110110001110100000111101001011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3927[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3927, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010010100110001111101000100000111011011010001011000110011010001101000111011111111111000001010100010011010110001000000110010000; 
out3928 = 128'b11101101000011101001111010000111001101100000100011110000011000101100111101011100110001001001111101000100110001011111111101110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3928[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3928, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100000101101111010110100010000100100111100000100111100010101011011011010001001101111010100010011101010010110110101011111111101; 
out3929 = 128'b10000101000000100111011001110000111110101100101111111001011110010111011100011110011001101101101111110110010100100001110100100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3929[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3929, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010011011101000100111111110101100111111111100111101100100000000011101100111000011000101000011000110111101011011100101011111; 
out3930 = 128'b01010001000010110001001100001110011111111110111001000010000010111111100011110010011011111111011001010001000000010010001001010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3930[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3930, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010011000110001010110110101111111010111110100011110001011010000000111001111110101010001000001000010011111000001011101011011; 
out3931 = 128'b01111000001000110000101101101101110110011000011100010011010010101001011010000100101011110010100000100011110110001101111000001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3931[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3931, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001111100000011000000000110100010100010101001011000111001101100110000110111010100110111111110100010000000111101000011111001100; 
out3932 = 128'b00110011000100001110001101100001011000111001101011011001001101111010111011101101001001101000010001111000110010000010010110111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3932[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3932, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110011010010101111100111010010110111000110101111010111000110100100111110110111110000000100000100111011101000010111011010110010; 
out3933 = 128'b01100001001100110100111101101010111100011111011000110111111011100101100011111101111101001001111110111110000111111111110001010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3933[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3933, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110010011100000100100101011101111110011100101111111001101011001000010100000100101101010100011101111101000001001111100100010; 
out3934 = 128'b10111101111111001011000111000111101010101010111001101010010110010001000110000100011011011111010001000110110100010010001100001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3934[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3934, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101101101011111101001111011011001111100100000000010100001001001011011110100000101100100000000100100110100001111000011000010101; 
out3935 = 128'b01000001011011111001111101001110110100110000001011001111000000011001100101000011101110100011111010000111011001011010101010011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3935[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3935, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101001010000001100111010110011010010011111010001101100110101010111110111000001000101110101111101100000010010001101111111000; 
out3936 = 128'b10000111111001011011000110010010111011111111101101001101010010100101001010011011110100010011101100010010001101001000001111011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3936[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3936, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011100000011101010000101011110010100000111110100000010110100010000100011010011110011101111000101101100010001010100000001000; 
out3937 = 128'b11111101011000111001011010010110000110111110011111101111011111011011100000100011000111010011101000010001010110100101101011000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3937[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3937, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010101110011011100101010111101010001001010101011011100001000101000001001110110000111011001011000111010001000011100011111010000; 
out3938 = 128'b11000011011110100110010111001101000001110101101011001010010110101110101110011011010111100011001101100011000111001111000110010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3938[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3938, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111010100000111010101011011100100101000011111101000001101000101000011110110011000100100100010111111000111101010110000100100; 
out3939 = 128'b00010110000011100001011001100000101111010101100111001100110010100101101011011010111001100100011111111100000000011110001111100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3939[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3939, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100000111000110010110110100110111110001101100110010011110101100100110011001001110000110100101110111110110011000010111011011; 
out3940 = 128'b01000011101010011001110011110010110110001000001001010010111110011010100010001000001001101101010100100100110001001110010111111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3940[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3940, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101101011111110101101000011110011100100100011111011111011111000011011101100000110001011000101111000001110010110101010000110; 
out3941 = 128'b01110111111000110000001111001100101011111011101011101011001110101001010111011011101010110110010110100001000011010001101110000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3941[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3941, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110001001111100111010010100010110000111110101000110001100100000001011001010111001010100101100100000101111000000000101010111; 
out3942 = 128'b00101000110000000001011001111000010101111111111010011101001100111011010001110110110010111101000111101001110111101111111111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3942[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3942, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100101111011001001000111010010010100010010111010110001010100001001101101010000011110011001110110011010001101101000110010011; 
out3943 = 128'b01000010001011000100101111001101101000101111010000001010011010001110000011011010000110100010110110111101110000100010101111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3943[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3943, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100110101011001101110001000010001101100111011101001111000111000101010000001100000100010000010011110001101010111010110111101; 
out3944 = 128'b10011000010111101111110100101101011111011110011110000100000001001110100111001000010101011000111010001000110010111011101111010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3944[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3944, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100010110011011010001110101111000110011010011101100110100110010010001111011011100111111100101101001000111011101001100010110; 
out3945 = 128'b11111111110100100001000001001100100011000010101000111011001110011100101100000100101111101111000011001110111111001110011100011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3945[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3945, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011000111000001001000001101011001100110101010011011011110111001011011101010001100111111010010011101011000100000011010000011; 
out3946 = 128'b11100011011010101101111110110010111111111111100100000101011011001011000001010101111001001010011100111111001111010100100001110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3946[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3946, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001000011001001110011010110011001111101000001100101111001010110011010000100100010100001010111111101110011000100111000110011; 
out3947 = 128'b11001100000111010001001000100001110110000110000000010111101111001111101000100000000000000010100101100101111000000010000001111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3947[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3947, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010100101110111011101010111001010010011000010011101011101100001011101011000111101001110111001010011100001110011011111001010; 
out3948 = 128'b01001011111110010001111000100000000001110111000011100101000100100111011000000111100000000100011111110101011100011011100100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3948[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3948, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111110000111101110000001101101101101001010111011111101000011111110010000001011110010011000101000011101100011010110001011001110; 
out3949 = 128'b00111110001010100010010011010110010000110010010001101001110111101111101000101111100000101000110010011001000111100110100101111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3949[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3949, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100010101100111000011111110010111001001111010111110111010001111000011011001001100000010010110000111111001010111011010001001; 
out3950 = 128'b10011101111010111100010101100111111101101111010010100111101000001100001011110001110000011110010001001111010101000010001000001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3950[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3950, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010011010110010000010111001101000101011100010011101010001001111000010111010111001101110111101010000110100101100010001100001001; 
out3951 = 128'b00011011111111010101101100111100110111001000001110010001100110010111001010110100011111100001010111100101001011111101111000110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3951[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3951, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111110100011110111011100111100101001101100111110001111000101110101110010010010101011100000100101010001010010010001010011110; 
out3952 = 128'b00000111100001000110101001100111000000100000111000001011111000000001101001100000111100001000001110000111011111000100101110110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3952[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3952, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101010011110011101101111001101000001010101010001101101101011000111001001011111011100100101110101110000001010101011011110110; 
out3953 = 128'b00011001011010111110001011010011100110000111101110101000111101111110011101001101110110101110111101111111010100111101010110111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3953[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3953, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111000011010001000110110110011110110011000000111100011010001110100010100111110111100101110010000001010010111110101111110101000; 
out3954 = 128'b00110110010000111010101001011111010111101100011010100011011000000000011000100010001010111000110100000100010111000001101000001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3954[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3954, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010111010001001110111100011111110110111101001100000011101001010101101101110111101101010101100001110100000110001110010010100; 
out3955 = 128'b11001010101110100100011011110010000011111001110010100100110101000000000101100000000000000011111100001100101000110010101110011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3955[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3955, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111011000101011100001011011100100011010101001011110010011110100011100111111010010000110010000001101111100111001011101011101011; 
out3956 = 128'b00111011010001000011000111010010000101111010001000000111100101000000111101101001011101100001100001101010110001010011010100110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3956[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3956, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100001001100110001100011110000010100000110111010000110001011100111110100000010010110010011001000111001100110011000100010001; 
out3957 = 128'b10101010000111101111011001111101101001100001000000111110011100010010001001110011001001111100001001101010111001111101111111110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3957[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3957, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110010111111100100001011001010110101110001101000101010110111100100110001000110100111001110101001100101110000110101100101100111; 
out3958 = 128'b01100110000111110101001010110100011000010100000101100110110100000101010111011111111100111111100100010010000111001101011001000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3958[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3958, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111001100100110001010001101000100011110100001000011101011101100101101001100110010010110010001111110101011010100101011110001; 
out3959 = 128'b11001011110001001000000110000110011111010001110000100001010011001010110101000011001100111001010011101100000100100101010111000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3959[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3959, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100011100010000111101100000101000011100101000100011001000100111101001010101110011100111100111001110101010110001010100010110; 
out3960 = 128'b01001011101011111000101000111001011100000100101101100000010000100101010001110111000101000110001100111011111110101111011111101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3960[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3960, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110111010000001000000011110100101000000110001010001011011110111011101110111001000001111001011111101110010001100011110111011100; 
out3961 = 128'b01110000111001111010010000010000110110000010100011111001101001001010001101100000010000000011010000100010000110011100110001111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3961[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3961, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101100000111100110001111110111100100011110110001011010100011010000101100111001101000100101001110011110101010011111101100000100; 
out3962 = 128'b01011000110001110010000011010001110101111011001111010111011100011100001111000110010001110110111110101111111100011010101010010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3962[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3962, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010001101101101010110100100010011011011000011001000000001110111011111001101000011101101101111000010100010011000001000000101; 
out3963 = 128'b01010000010010101011001000000010010110101111001001110110010001111101111011011111101111001010010111111101000110000001010100100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3963[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3963, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100010111010100110111101101111111011111101111111110011010001101001101110010001001001001000000010000111001011100001101011011; 
out3964 = 128'b10110100000001111001000111010011001001001111000101011000111110001001000101100011000010110000111100100100111010110111101010101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3964[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3964, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111110010110011000101001101111111001100110010101110100110011111101101110010011001010000010111000101010100100111101010000001111; 
out3965 = 128'b01100111000000100010101010111111011101011111100101001110000001101010001111011111011101110000100001000001010000000111010101101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3965[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3965, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010111110100000100110010010011101001000000010010111000100100010011111010110110011100111000101100110100100011010001101011100000; 
out3966 = 128'b01000110110100110111111110110000000011000010101100111100010010110011110111010101001100101000101000001000100001111000100010000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3966[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3966, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000011001111101011011000001000100100001001110101000101101011101110000101011100100101011000111101110001101001010100110111000101; 
out3967 = 128'b00000100010010011111001110100101110000000100011010111111101010011100111010100101000110110010011000101011111001000000011011010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3967[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3967, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001011101010010111000101010010100000011000001111101010101000011111110010100100111100001110011101110010011010001000110101101110; 
out3968 = 128'b10011011010011101010001011010010010101000101100111111011010011010001111111000011010101011111111110001011100000000110110111111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3968[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3968, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100100100011011100110000010001110000110001001101100101000100001010001111101101010110111000000010110100011100111011001001000111; 
out3969 = 128'b00000010100000110100101101001011100111110010100111011110000100111001010011101100110000001100111011100001010101011101100111110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3969[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3969, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000001000010010010110110111110111011000111100001100001110110011111100011001010110100011111111001001100101011001000010110100; 
out3970 = 128'b10010111111010100101111010001001100011010010010101000110110010101010101010100001110011010000101110010010111101011000010011000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3970[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3970, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000001010111100111000111101001100010110001010100010100101100010100100000000011100100000001010101010100000010000011001101111; 
out3971 = 128'b11011000100100001000100110001010001110000101110101110111101101101001011001011000101101000010011011100000101101100011010010100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3971[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3971, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011011100110000110101100111000010011101100101100110011001111111010001011110101100000001011011000100001111001001010101001100; 
out3972 = 128'b11010001111100100010100011001001101110001000101111111111111001111111101111110101111000111110101011001001010010000001000011010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3972[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3972, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101100101000101010011111001011100001100000110010100010011000011001000110111001001100111101110101011110011010000100110010011; 
out3973 = 128'b01100001111111001101001101101100101100110101011001010110010100010101100111011101011111011100010001000000010110111001011010101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3973[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3973, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001100000011000100110110101100001000011001111010000110011010110011011011011011101000111000110011000011000110110011111101010; 
out3974 = 128'b11101001111100110101011111010101100101110000001010101011011101111110110011010111101001100000001100111111000011111000001110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3974[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3974, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100100010010100010011111001100011010111010111110101001011001011000000110100110010000011110010100010001110000100000011111001; 
out3975 = 128'b01001011010010010011011100001111001001110100001011000100001010111010101100111101000100101110011000000100100001010000100011100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3975[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3975, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101011000100010110101010101110000101110000011000110111100110101010011100011110110010100101010010001011001101100100111000100; 
out3976 = 128'b11001110000100100001110011110110100011100100001111000011111001100000010010111000100110100001010010010111110111101010000100110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3976[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3976, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100111011100010001010000001101110110011000110010111111010011000101001110111100000001111010001111010100111100110101100000011; 
out3977 = 128'b11011001111011010110111010010010001010001011000111100100100111100101100010010011000010111000011111000100001111010000100001001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3977[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3977, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010100110100010110110100111101001011011000011010100110000100101110000010001010001100011111111000111011001101010100110000001; 
out3978 = 128'b10100010010000001101001011110011111010010001001100100111100110101010011101100110010111111101111011111100111101010010001110101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3978[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3978, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011101100101100001010110010000000101000100100010101111000101000010011010101010000010110111101100010000010001100110001001110011; 
out3979 = 128'b00000110000010110110011001001100100011010111010001001111111101110010010001100011011010001101100110100110001100101011100111001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3979[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3979, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101111101000111100011100000010001111000000011110100011011000000111011101001111111101110110011001010010010110010111111100100; 
out3980 = 128'b10010000011111100101010010011100010011001101101100001001001010010101101000100011110000001010001011000100111101101101101001111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3980[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3980, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011011100010101111011001111101010101010111110001110111111101101101111001011110001101110001000001111000001100110101111010111; 
out3981 = 128'b01010011000011010110100000101101010001100100110010001001001101011001001110111111001100111101010111101101101110100101100000111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3981[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3981, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001000111100111101110010010000100101001001011010001111001101101100100011100001010101010100010111111110011111000111000000000; 
out3982 = 128'b10111010101110111010101001000101111100001010011001101101110100001110010000000001100100101101100011001011100110011110000111101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3982[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3982, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010001101111010101110111100010011011000010011101111101001111101010000100111110100101000111101110101110101101001011101001000010; 
out3983 = 128'b11001010000111101001001100100110111111011111101110011100101110110110011010000100100110011110110110011101011011011101111110100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3983[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3983, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111010110101001101111101101101111111011001101000100001001010010100100111111000101100110101010001101101111111100111101000101000; 
out3984 = 128'b00101001111100000010011110100000100001111000111110011101111000101000011110000100000001111101010011011000110110001111010011101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3984[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3984, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001100110110101100011011101100001001010100000000111001100000111001001011110100011101111101111110111001101010000000101000011; 
out3985 = 128'b01000110001001111010101001000111110000001000100001111001100001001010110101010110011000111001110100000010010111010101001001011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3985[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3985, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101000110111110101011111010010011111101110010111001101000010001001000000011011001111100111111100100110110100110111111000101; 
out3986 = 128'b11111011101001111111011010010011000110111111000111100001010010001101101011110010000001111010001110100010110101110000101110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3986[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3986, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000111000011000001000111111010101100101110101111111100011111100011011000101011001011010011000111001000000001010001000100101; 
out3987 = 128'b01111000011100111100010100110001001100011111111001101110000101001100000000100110011000011001001010110111101001100101111010010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3987[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3987, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111011011101101111011001111011101110110100101110010100010110111100100111101001111000110111101110100110100101100001101010111; 
out3988 = 128'b00000111110110010111111100010100011001101100011010100011100000011100001100110100000011010111000100101001011010001110001010110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3988[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3988, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010010000010110101110101000001101100000111100001111010110101011000011010000101010100010000110010111111011101110100111010111; 
out3989 = 128'b00000010100101110001000011110000001010100011010011010110100111100110011101100010011101000100111000001101110101110111110010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3989[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3989, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100001110010001100101110111000100100010011001101011101100000010000011011010011101101001001001110110100010000010101111100101100; 
out3990 = 128'b11000110001111110001101110001000011101100000101101101101110001010101100100001110011001110110000010001111001011010011001011100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3990[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3990, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100110010111001111101110000010101100111100000011110110010100000010001001100000001000000001100100111100011100111011001111101; 
out3991 = 128'b10011101011110111011111110000111000001100111110110111000100110100110010111101010010101011110010000010101011110100011011000000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3991[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3991, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000111111011011111010011000110101000001010000100111000100101110110100101101000001111011001011101110001110010111111000001101; 
out3992 = 128'b00011110100111010011101100010110001011001001100011101110000101001101101011110010011000101001011101010101001110011000011101010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3992[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3992, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100101001101110101110011010101101110011100101110101110010111001101101111111111101100100011101101101111100000101100101111011; 
out3993 = 128'b00101010110100100110000011110000111001000110010011011110111101100110000011010000010001010110000100101111001011010110011101110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3993[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3993, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000000110000110111001101111100000100001111010001111101001001101101100010101100101001100000111000110111001000101110010111001; 
out3994 = 128'b11100101110100110110100100100101100010011000110011110000000101100101001000001101000000100011101110011000000010011111010101111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3994[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3994, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100000100110111000000010000101110100101011001001010100011111111000011100101101101011100110101111000100111110010001011111100010; 
out3995 = 128'b00101100100110001100110001010111110001110111000110100010010110010101010001011110010110101101001000111111101101001101101111001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3995[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3995, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010010101011100001001111100001011000000101111010001111110100000000111000001011000111111110011111101111100110111000000110110101; 
out3996 = 128'b10101100001111100010101011111110100010111000001100110010010100010101010010100011100001100101010100100000001011101100000001100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3996[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3996, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111000100001001101001101101110111100011001100010100010111100110011001111011000000111011010111100011001111101000001100100001; 
out3997 = 128'b01101011111000110111000001111111011100111010011111101101001100001110100001111101101000001011110111001101001010000010001010101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3997[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3997, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000110101000101111000111111011110101110101001101111011000001101100000011000100111001010100011000010010100111011000000111101; 
out3998 = 128'b01101010100111110001101100111010001011100110100000100001111111100011000010101111001110000010110010100111111011000101000101100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3998[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3998, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111011010010010010111001111101001100010100001100111001000110011001101100010011110001111111010101011010011100110100011111011; 
out3999 = 128'b01100011011011010100011100111001111111111000110110000111000111101000011011110000110001000110011010101001101110111000101101110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out3999[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out3999, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010010100000011001000111101111111111110110000111111001000101110000100001101101101001010010101001000001000001011100001010111; 
out4000 = 128'b00010010011100010100101011111000000101000011101100010110001001101101011001010111111111111100101101110000010001111111001101111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4000[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4000, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110001110100011110101110100000100001101110011010000010000111010011001100011110000000001001000010011010100010011111001101001; 
out4001 = 128'b01001010101100100001000010000011000101100110011101000010110101011011011010100000011011111001011010100001100010000001011010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4001[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4001, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000111001100110010010011001000110100011111010110111000101000000000101000010001010000110011111000001001110110100101110100000; 
out4002 = 128'b01101010101111111011010111001010110010011101000101110011110001111101010101100111000111111001100010011110011110000000110110000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4002[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4002, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011101001000001110110110001011111011010001000110001001111000010100010100111001110100011011101011101111011001001110010110111; 
out4003 = 128'b01011100100100000101111011000011011000011001110110100110101011011000110000101001111011000101001110110011011000001101111011001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4003[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4003, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011011100001010011011010101000110000111100110010001010110110000011100100010011111011011110110011011000110010110001111000110; 
out4004 = 128'b01011010100010010110001010010110010010000101011111010010011011111110011101100000010110101001010001001110110010110011001110010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4004[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4004, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110111011000010100111111001001000011101000111110100000111010110000010010010001000011101110110101101010110010001000010101100; 
out4005 = 128'b10010011100010011000101011000000100101111011111010111100100101110001001000111111111100100011100101011110101010011100010010101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4005[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4005, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110010000011100001001001010101100000100110100111110010110000100011011110000011000111110010001000000000110110001101001100011; 
out4006 = 128'b11110100000010110010010001000110000111101100110111101011101101011000111100001001001100001101100100000100000110000011011000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4006[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4006, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101001001110001001000110010100011110011101101010111111111001111100011111111011001001010011000011100111010110101001011001011001; 
out4007 = 128'b10100100110101010100010010111000110010111000101100010001001010011111001110111010011011000011101111110110101101011000101010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4007[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4007, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111100001010101011000100101101001000000100011110101010000101010011110110110000100111111010000111110101001101010101011111110101; 
out4008 = 128'b00111111011101110010101000000100110001110111111000000011001000010001101110101010010110010000101110111101001011100010001111000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4008[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4008, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001010110110101100111110111101011111101110110110100110101000110001101011110000111110001110101111010001010011101000100110100; 
out4009 = 128'b01101011100001101001001100000011111001000101000000110000111101000100011101111100111001011100111010001101011001100010000101011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4009[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4009, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010011111000010001100001001101001001010010001101101110101110110001100001111001000100011111101001100001011000010100101110101; 
out4010 = 128'b01101000000010110111110001101000100000101100101101011010101000011000100000000101001110111000111111001000010010111001101000111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4010[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4010, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111111011000101011110111110010101001111011111101000010000010111100111100101110100110110111111110101000001100000101000000111; 
out4011 = 128'b11001010110100010100001000001101100011011100110101010101110001011000001111100100101100001011011100000000110111010010100000111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4011[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4011, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100000000101110000010011110101101110000000100010110101011011111100100011011010001001011001101001100000001001100000011110011; 
out4012 = 128'b00010011011011110010110111101000100111010001011010001010010011111111011001001100100101101000000001010010010110111111100111110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4012[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4012, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000011011010101010100101111010011111000110000100011100001100000110101011001011011101110001011110101011100001001011000100101; 
out4013 = 128'b00100000001101000110010010101111101011001101001101010111011111010000100110001011100101000111011111011011001001011100010010110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4013[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4013, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001001001001011100000000110111001000111111111000010100101111011001001011011000001101100011011111111110000101010100011011111; 
out4014 = 128'b00011011010011110011110000100000110000010110100101011011011000001011110110110011000100011110110110011100101010100111111111000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4014[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4014, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111101100011110100111010110111100011001110010110101100000110010100011100000100101010011000010011100011010101000000011111111; 
out4015 = 128'b01101100100101000111100000101001001001111010111101110101100100100101010101011010000110001110101000001011010000010001110011001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4015[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4015, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010001000010000000001111010100001100111010010010100001100110010000010011010111100010001100000110001110100000100111001011100010; 
out4016 = 128'b11101010111110011101011010001000010111010100010110011010100100110011101001000001110000011111110000101101111100111010011100101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4016[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4016, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010010011001101100111010010111111011111010001001011111000000111001011111000001101000110111010001100100101100101010010001101100; 
out4017 = 128'b11101110101110000001010001011001111000111101110100100111101110111011010100110011111010100111010100000110011011010101111111111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4017[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4017, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101000010010011100001110100010111111010101011101101010011110000111010100111100100001000101000011101110100100000111000111000101; 
out4018 = 128'b10011110011101011000001111111011110010100100110101010010010100000110010010101100101010101001111100001010101010110001110011111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4018[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4018, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110000110110001101011010111100001101011000011110111000111001111001101101110011111110001110000010011001000111110010000100011; 
out4019 = 128'b11010111100001101011111001101101001011110001010010011111100111111010111111101110011011101010110001000001111100100001001011001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4019[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4019, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000110001011100010001111101011010100000100111111001110001110111001011101010011101010000011010010000110100010101000111100000; 
out4020 = 128'b01101100101001111001111111000110010011011111100011001110011001010011111000011101111111010000110010001010101111000101101000110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4020[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4020, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000011001101100111100000100011000001101110000111100010001011011111010011111110100101101010010110011010011100100110110101110; 
out4021 = 128'b00010010101000010111010011111100101100010000010000001110111000111011001111001000101001100000000111010011000010100100001000000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4021[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4021, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000010110100101111110100110010000101011010101000111111011111000101100011101010000010000010010000001110110101010010000101110; 
out4022 = 128'b11001111111100101111111111111100101010110100100100101110001100001000110010010010111001000111111010111100110101110101010010000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4022[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4022, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011001010011110001111100000111111110011010001010010011001010100110111101111100100111001001100010001010000110101110100001010111; 
out4023 = 128'b10000110100010011011101000000111010000111111111111010001110111110100000010011100010000010111101111110000010100011011011110011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4023[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4023, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000010110111100010011100011011011101000110111010110111011100011101001110110000100001001110101010011111100110010011000000111; 
out4024 = 128'b11111010011110101110011000000100000110100110001001100100001010101011000110101110111011101101011100101000111110110000001111001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4024[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4024, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001101101111000111101010100111100010001111010111110011100001011100100101111011011010011000011111011110100101001001111000111000; 
out4025 = 128'b01010100101100100111101101011010000001010010110111100101001000110000100111100111001101110111001100101000110010100101101000011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4025[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4025, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001100010010101100100111110011110001101000110101011111100000001110000111000000000000100110110101100001100111010010000111101001; 
out4026 = 128'b10001110111001001111011010001010101110111101001111110111010000011110000100010011011111110110001110100110111110100010101001011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4026[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4026, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111001101110000001011011001001011101000101010111011011101101010001000001101100110011011110110011010110011100101000010000010111; 
out4027 = 128'b00000000111001011001111000010000011000110100001010100111110110000101010001010010010010001111111010100110001011110101100011010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4027[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4027, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001110001010000111101001010110010011001100110100000001111001001011011100000011111111111010100001010001111010011001101100011110; 
out4028 = 128'b00110101100110011111111011010011011010010100101010110000101110011101101101010000011010100101001101010001111110011010001100000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4028[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4028, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000000100110110001100011111101100000010111111111010101110010011100011110011110010001111001110111010110111111010110110001000; 
out4029 = 128'b01101101111000011000000001111000001010011011110111101011000111000110011010011110011010011000011111011000000000100110000011100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4029[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4029, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111101001100111101101001101100011010011110111111100000100100111011111100111111001011000110110110001111100011111011110101001; 
out4030 = 128'b10111010001100111110001001101101000110000101100110111000100100111001010001000010110010000011010111011000010000100000100111100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4030[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4030, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110000010110010000101001011010101100010111011000011000001101101011101111001100001011111010000000110010110111001110100010110; 
out4031 = 128'b11101111010010111100110010011011100000111101100111110001001111000100100010011101000000101000100111100100100101011010000100101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4031[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4031, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001110110100101001100001111010111011101010011110000111011110011100010001100001011101000001100010110110100100000010111011101111; 
out4032 = 128'b00101110101010010011100100100010010100010101001001101101011111101000100011000000001100110101111011110101111001101001111010010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4032[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4032, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111100011111100101010010111011110101011010000010101011110101110011101010100001110010100100011000111011010100101100110001110; 
out4033 = 128'b11000100000010111110000110000110110100001000110001111110011011010011010111101110101101110111001010011001101001111011010101010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4033[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4033, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110100001101100000101111011001111000010100000110011101110011011001011100001110111010101111001100000100010100110011010010011; 
out4034 = 128'b10001100100001101100110100111000010001111100000001101001000000000101010100010001110101010110111100100001110111101010100011100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4034[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4034, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011100111010111110111010010110110010010000100010110111001101111000000000111010110000001100100011101001000110001111110110010; 
out4035 = 128'b11000111101010011001010101000100011010110111000010111011100011000000111110011111011101001000100010001110010000001110011100110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4035[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4035, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110110000010111100111110100111110111110100101001011000111000111001011101100110100111000000100011100011011110100001010100001; 
out4036 = 128'b11101100111010010101001001011010101111000011111010111001001001000000111000011100001110100111111011011010111011101111001000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4036[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4036, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100001001000100101110101110010110110001101100111000111111111110011010110100011010000111000101100011010111110101110101100011; 
out4037 = 128'b10111111111111010110010011000010011010101101001011011101110010010000111011010001100010001010100010010000011001000111011000110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4037[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4037, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000001111001111110101001110010000110001100001100111010000011010001011010011011101110000111000000101001101110010111100101111; 
out4038 = 128'b01010101000110000110001111101101000001011011011001111000001010111001011100111010110110111111001100110001101011101000000011111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4038[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4038, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110111110011001011010111110011010001100110011011011011011001001001110111111010000000010010101111110111010110010110110101001; 
out4039 = 128'b10011011110001100010001100011101011110011010011101011010001010001000101000111011101011000101000001011001001111000010001001111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4039[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4039, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010000010100101110111111011001011001100000011100100101100010011111001010010101000111000011100001010110000000011100010000000; 
out4040 = 128'b01110010010110001011000101011110101101011100001100000010011010001101010001100101111000001010100100011111110111010110010111110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4040[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4040, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000101010111110111111110000111010100010110011011111110111101001110011101101111000011100000000111110011000000001101100010010001; 
out4041 = 128'b11001110011010110111010100110001110010001001101110011010001000001110110101110000010110101001111110110111111111100001000000111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4041[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4041, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111010000100010010101100000101011011011110001001100010000000110100011110000100010100100100011011001010101000001011101111101; 
out4042 = 128'b11001001001010111101110010110000001001011101010111011101111011010111000101000111011000011110001000111101001000110001000011111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4042[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4042, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101011101111101111010010111001001100001111010100100101011110101000010011011110110101110100011110001001101101101111011011010010; 
out4043 = 128'b10000010100010011110011010001000011000101010011111001010101000001100011010100101010101001101010000010001010000011010101100001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4043[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4043, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100000111100001110100001110101011110010110011110001101110101100011100000110110001000101000100010010001001100011010010001101; 
out4044 = 128'b10010100111100001110001000101001100111000101101111001001010000001011011010011010001101000110100000100001010110110110100100000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4044[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4044, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100001111011101111010111110001001101100000110011001001010111100010111011000011000110110000011101101011010111101011010010111111; 
out4045 = 128'b10011011111000011110010011000111010111101000100100011010111010000000011111100011010100100101000000011111010101001100100001110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4045[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4045, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110110010100111011101000000010001011010011110001001001110011010011000010010001000110100000000001101101111111110100100100001000; 
out4046 = 128'b10111011001001111111011100110111101001111000000101011110100111100111100000110000001000100101000000010000011011001010000010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4046[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4046, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000001010111010110000100000100010111011111111100111011000101101000011100001011001101010011010011011110010011000101100000000; 
out4047 = 128'b10101011011000110011010000001110010010101100101110000100000110100000010010011011010011001010101010001010001100100111101110110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4047[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4047, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000101100010011000010000111011110000101100001101011010100001001000110110000001100001011001110011011101011100000011111101101100; 
out4048 = 128'b01101100101010101110000010111000011000111100001011000000101100001001011100110100011010011001001011000011101100110011010001011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4048[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4048, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110011010011011000011000000110100001010001110010100001111011111011001101110001101000100100111101010010101010001100001010011101; 
out4049 = 128'b01010110100100010110100000000101111011111110110011110000011101100000001011001110000000111010001001001011110101010000000001010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4049[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4049, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111111000100010010110001100001010011101011111000100010000010000101110101010000000110100000100111111110100000000111011111110; 
out4050 = 128'b11111100011000100110011111011110010111100010111100011000101001000011010011001110010001011101000110100101000111111000111001000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4050[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4050, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111110011100011011110010100011101000010100010011110101110100001011010011000111011100001010010100100110010011111001101110010010; 
out4051 = 128'b00000111010001011011010010010110101000000100100111110001100010110110111111000011110100010110110011000101010100100101110101110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4051[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4051, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001101100110011000010011010111110000110100110000110101011110011110000011101000110111111011010100000100111011010011011100100; 
out4052 = 128'b01010101110001011101001101101101010001101000001100010110001100100110110101011010100100010100011011011101010010101111011010010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4052[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4052, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010100110011000000011010011001101101110100100001011001001101100001101010011100101000110100000011010001011010000111011101010100; 
out4053 = 128'b01011011000110110000001011110111100011100001010110100111011000001010011110100000111010011110111100010011001000100100100100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4053[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4053, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101101000010111010000010100101110111010110001101000001000000101010110000010000110110010101101101000111001000101010101110000; 
out4054 = 128'b11001011011010110110110010101010001010100110011010000100110100011111001011111010111011110001110101110100100101001010000100001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4054[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4054, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100000011001000100000101110011011010011101111101110111010000010001110010101111011010010010011101011110011111011011100111110101; 
out4055 = 128'b11110001101111110010101011001010001010010000001111011100011110010101101111010000101100101010100001010011001011000001010010110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4055[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4055, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111100001110111000010111010110110010010010010000000100001111011110000110110111110000011000000000101010101111111101000000100110; 
out4056 = 128'b10110000111010001000001100010100011001110100110110000101001110110000101110111101100011001010010001011100110001010011110010011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4056[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4056, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010001010011100101000110101100000011110110001010010100101111101110000100100010100010010001101000110010100010100011000101000000; 
out4057 = 128'b00010001101111001000110100100100001001001000100011010100111000101001001110101000010000110110111101000001100011001101111100011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4057[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4057, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000101010100001010001111000110111111100110010011001110011101111101010011001000110110111111000010001100010000101111111111100000; 
out4058 = 128'b00111101000011001010110100010000010010111001100110101101101010110110111001110110101001011111001100000001011000100111010000010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4058[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4058, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100001101010001101000100100100011000011110001100001111110100011010110001001011100101100010010001100011010100010001100000100; 
out4059 = 128'b01001100100001111100001101000100010110111111010110100001001111000100111100110000111010000111010101011000111100010111001000010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4059[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4059, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111100111001101110011100010111111000000110110001101110101000001100101100111100100111010011100010111111100010011111010100100; 
out4060 = 128'b01111111110011011101000110100000001000110010101101000111011011001010011110011111100000010101001001111100001110110100111111100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4060[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4060, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101011011000101111001110111101111100011110100001110110111001110111101100001111110100101111011011111110010100100001100011000; 
out4061 = 128'b01001000110001011000111101001000110110001010100101010011000101000100101011100110111001000011000001100000011001011100010101110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4061[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4061, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111111000100100101100010000010001011101101111100010001001000010110011110010111001001011000000100000111000001101010100001001; 
out4062 = 128'b00101100010100001000000110010111010111001010000001000100000011000000101000011001001101100011110110101111000011100101101001101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4062[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4062, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000111111101011111110001011010100011001101100011101110011010000101011100110100000000101110010011000110100011001001001100110; 
out4063 = 128'b10010101101111101011101000101011011110000111101111011010100100011001110001111111111001101100101110110001101011010011111001111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4063[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4063, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011100110111100110101100000101100101011010110101001110010111000000001110000111011010001011110101011010001101111010111001011101; 
out4064 = 128'b11101000101100111110101100111110111001011110000010100011011000101010000110000100010000011010110101100100011100001011000011100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4064[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4064, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110100011101111100110011011100100000000011100100011001111111001110010011111101111110010110011011110000110100010100111100011011; 
out4065 = 128'b11001111101111101110100101111001011001011110010100110001100001001010000100010001000100101001110001111100100011111011110111101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4065[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4065, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111111101110110111110010110111001110000001001001010010000111100101111100001110000101001010011011000001100011100010000111011; 
out4066 = 128'b11101101011001001000011011000001001100011000010101101110101010011000011101100110011010001011001010010100111001011100000111100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4066[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4066, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001010110000011010110110110100010011100001100111101000000111110110110011100000100001111101110101110111111100011011011001101; 
out4067 = 128'b01001011001011110111010101011101111001000111100100101001110011011001010111110011110000000011100101111011001010100001100010111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4067[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4067, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100100101011001001101011000110101010010001011011101110110011101110000101001010010110111010000111011011000100110000000011010; 
out4068 = 128'b01100101001010001100110000010001010111000000010111011100111000101011010001011011111100010111110111110100001110100000010101010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4068[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4068, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001101100100011001000100011000110111101100010110011100000100110110100011111011111010010101110010001110010000111111011100011; 
out4069 = 128'b01101001010011011111001011100001111001011010100111000011000000000000110000000100001011111000010001110001011001001101100010011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4069[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4069, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110111110111000111001011100001001000001011001111001111111001110001000010101011001111001000001101000100011000100001000010000; 
out4070 = 128'b10101101011011111110100110111000111111110011111010101110110101011100111001001101110010100000110111111011000010101111011001101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4070[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4070, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101001111001100110000000011011001100001110011111010110001101011100101100011100011110110000111010100011010011000111000110100001; 
out4071 = 128'b00010100101111011101100100001111100000100001111111000000101100010101010000111110111000001100010100101111011010001101001110011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4071[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4071, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110100000000100001101001011100111000111001111110011000101001010001110100110101000101000111010011010110011100101111101101100; 
out4072 = 128'b00100001000100011100101000011101000100111101111001101011100111010111111010111110001101010010010001000100110100001110011101001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4072[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4072, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110010100011010011100010110101000001010100010011111010111011110101101110010001101011000000000100100011000100000000010011110; 
out4073 = 128'b11000100010011100100000111110100001100111110001111110111010011011110001011111111101101001001100101011000110011100001111111111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4073[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4073, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101000100110110100111110000010001000101101000001110111101111011100001010001110000100110001010111110110111111110001110110111001; 
out4074 = 128'b11010110011111111110100000001001101101011001110000100000111111110101110110110111001011001000111001010000000001100101100111001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4074[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4074, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001000011100010111101101101111011111011001010011111110011101010010100101000101100011111000000110011100101100000110000000011010; 
out4075 = 128'b01001011001101011000000011111101001111100111101110101111011110101101101011000110111110001010100110111110111101001110111101101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4075[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4075, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001100000000101100001100110100110111011010101111000011111001001010010010000001001101110101001101101011011111100001010000000100; 
out4076 = 128'b01100011101000011010011011001000001110011000100101110001111101100101001110101010000011110000101001111111101010010011100010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4076[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4076, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100000100101000101001101100111011100100010111110010011101110100010110101001110011010010111000101010010001001100001010010100010; 
out4077 = 128'b00110011010011110100110111111001000010011011000110110111001110110110001010100110101010011011111111011110100110100001110011010110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4077[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4077, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011100000000101011011010000000011001010001010010000001000010010010001111100001101110001000001101000001011011110000001011100; 
out4078 = 128'b00001010011110011111000111000010001001011000101000110111001011110001110101100001001100010111011010100000001001101001100011010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4078[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4078, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010011111100110011100110010101111011111001000101101001100110111001111011010100011011111011000101011101001011100000101010111; 
out4079 = 128'b01100010111110001110010011110010011011100110111100011011000011101100101100011011111000110001101000010111101101010011111111000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4079[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4079, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110000110000000001100001101000110100010011101001011001101001110011110101111001100110110011000101111010110110110011001101010; 
out4080 = 128'b10110100011010011001000010001011100011101001011100100001101111000111101001100001101001000100111011101010001010101000111010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4080[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4080, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011101001101101001100110100100100001100100100101000010110010010000000101000010011111100111111101011100011011100000001010111; 
out4081 = 128'b01010100101010100100111011001100000101001001111110010001000101101111101111110010000011001010110100010010100010010111110000010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4081[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4081, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000100001111011000011101111001110001100111000010110110111011101010011100100000011011110101000110100010010001111010011101010110; 
out4082 = 128'b01101101100000011010110101011011111101001101000010100010101010100100001000000011110010111010011110110001011110010001100010101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4082[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4082, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011101001010001110010000000001110110010101101101110100100101101101001100101110001101011010110111011101110100010000011011000111; 
out4083 = 128'b10110110001011001001110111110100111010101011011111010011110011110100000110111101001100111010000110100111000001001000000000110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4083[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4083, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110100111011101010101001110110111001011001111000011010111101110101000000111100110001100010110111101110011001110110101011010; 
out4084 = 128'b00010010011100101001110001010001101010101001011111100110100011100000000100001110011000110000011010111010100100000101010101100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4084[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4084, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111101010010010011010001011001100110011101010000000011111001101100100011111110111110101111000001110111010110110101001001010101; 
out4085 = 128'b00001100101101110001110110000001011010010010001000101000000101101011101011010001000111101001010010100010000101101000011111111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4085[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4085, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011001110001111001111001001111110010100110100010100101111011101001010010000111010101100111101100100010010100011101111100101101; 
out4086 = 128'b10110111011111010001001110001101100001110101010010011000000101011010000000001101010101001101100100000111000010111010000110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4086[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4086, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111100100111110111010111101001110110100010101110101110101110100101101100101010101000011011101010010000010001100101011100001; 
out4087 = 128'b11101100100000110001011100101101001110111001110100001110000011010000111110011000111010001100001001011001101100111110100101111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4087[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4087, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000100110110001100001101001011001000100001001100101001000110111100010000011111101111011001011111100100110010110111001011000; 
out4088 = 128'b01011100100010110110011111100100101110011011001000011110001101001111010000000111000000100000000001110111110101111011010010110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4088[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4088, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011111101101111110111000010010101100010011001110110111101000000010000010100010100011100100010110111010110111100011011110011100; 
out4089 = 128'b10000101010110011010000101000101000111010101111001001011011110101010011010100001101110110010101111110110001011111110111101000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4089[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4089, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000101000010000100000100000111110001100100001101011110100010100111110100001110001100001011010010011011001000100011000100011; 
out4090 = 128'b00101001101100010101010001010111100000000011001011010000101110000111100010111111111110001001001010011101001100100010100010011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4090[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4090, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111001000101111011110011111001110111001101000110110100100101100111110000101001010010001101000101100100010100100100101100001; 
out4091 = 128'b10011001010001100000100101001010010010011000100000111111001100010001110100101100000011001111110101111100111101101101100111001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4091[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4091, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111111010000000111100100000001100010101100001110111101000101001001110010010000011000010011100010001000010100111000000001100; 
out4092 = 128'b11111111111111111111110011001101101110111011110010011000010000110111101100000000110010001010000111000100011101011011110000111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4092[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4092, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001100111101110000111001000100001010110111010110000000010101011011001001001100000011011000010100111001110001100011011010011010; 
out4093 = 128'b00000111011111111000111111010011100000000110101100111101000101000010100010111100000110010000101010010001101111000111110000111101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4093[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4093, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110011001011001100101110000110100011010001011101001011110100010101011011110000100001010000001000100111010100010101010101101; 
out4094 = 128'b01110000000101001111100010011110111110111011111111100011010000000100111100001011101110111110000110010001000000010011001011110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4094[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4094, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101000001011111010010011000010011010001010100100111001110111101011001000100100101001000110011100100010001000001000000011011; 
out4095 = 128'b00100111110111110011001111110001001110110110110010010000011011000010000101011001000010111001110001011101001000101100011010011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4095[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4095, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111101100100011000100001101111101110101011100111101001110001011110010000000001110001101100001001010001000100111101111100010101; 
out4096 = 128'b00000001000011110001000111000001101000011001011111101011000010011010001101011001011101010011111011001000101011101101011101100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4096[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4096, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010000110111110010101010001110000011110000000111110101110101111111000001101000011000111011110001111111010010100010110011000; 
out4097 = 128'b11111001101110101110000101000010110110001000101011001111010110110111111111001011111001010101101100100010101111110110111010010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4097[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4097, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111; 
out4098 = 128'b10001010111100101000011000000001010000101111011110000110111101000000100100110000011111000001101000111111011111101010101010101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4098[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4098, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000111001001111000100010000010100101110100011100100100001000010000000001001000100001000000000100000010001000001001011001000; 
out4099 = 128'b11111011010001001011000100111011000111011111000100100101101101011000101001100110001010001111001101011010010111000110110100011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4099[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4099, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110000100110000010001101100000011010000000100010010000110001101001001110110011001110010010011001111001100011110000000100011; 
out4100 = 128'b11010011011100011111000001011101000010111011111000110101001110110001111011100100101100011101111111001110011011001111101111001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4100[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4100, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111111111011110111110101001010110111010001101010010100010110001101011110011111000100011111001010001000010101000000101001111; 
out4101 = 128'b10011111101110011000101001001010110010000010001011000110010010001001101100010110010011110111110100111011000011001001011001010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4101[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4101, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111111110111101111101010010101101110100011010100101000101100011010111100111110001000111110010100010000101010000001010011110; 
out4102 = 128'b01100110001100010101001100010010010101111011111100000010000011101000100100011010011110101110101010010101101100001000000111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4102[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4102, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101111011000101101111110100101011110110110101110100100101101001010111000010100001001000111011001011110000110100000010100101; 
out4103 = 128'b10010110110100001001101110011110100101000101110011101100010001011100011101100101010000010101000000010101011101001111101101100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4103[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4103, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011110110001011011111101001010111101101101011101001001011010010101110000101000010010001110110010111100001101000000101001011; 
out4104 = 128'b01011001100011111111110110001010011100111110001101101010100101000111110010010011101001000000111110111100001100001110011101100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4104[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4104, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101101010101000101010000011011111000101010111101100111000001010100100000111000111100100110010100000111001000100011100001110; 
out4105 = 128'b00111111111011001100101111110001111101000011111000011110101101100111100111000000001011101000000110010110001000010110111100010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4105[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4105, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011010101010001010100000110111110001010101111011001110000010101001000001110001111001001100101000001110010001000111000011100; 
out4106 = 128'b11111001001101011011100001001001001110111010111110011000011011100100000001001111111111000001101010101011010000100001010100101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4106[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4106, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110101010100010101000001101111100010101011110110011100000101010010000011100011110010011001010000011100100010001110000111001; 
out4107 = 128'b01011010111111011001110101010010111101000101011100010100011011111101111000010010000111100100111011000000010101000011000000110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4107[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4107, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111010011111011000101001010001000110100111101011001101111111011011000110101111111100001001010001000110010110111110111101010; 
out4108 = 128'b10111011100010100110010111011011111110101001100111101001111110001101000111101111001000110010001111000111100011011111001111010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4108[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4108, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100100001001000011111000101100001110111111010001101110001011001001001100110111100000101001010011110011111111011111001001100; 
out4109 = 128'b01001011000001100011010100101100110111010010111110010001110110011101100010000100001011000111000010110101110010010001110010011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4109[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4109, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001000010010000111110001011000011101111110100011011100010110010010011001101111000001010010100111100111111110111110010011000; 
out4110 = 128'b10100000001111000110101001101101100001001111101100010011010100010010011010000111001101001000001001111010111110100011111011000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4110[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4110, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000000010011111101001000111110111000001101000001001101011001011011110010110110011010011110111110110000101111011110010101000; 
out4111 = 128'b10110011011100000100110110001101100110101000010111010101110111011001011100011000111110111010111011101111101000011001110100000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4111[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4111, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010000000100111111010010001111101110000011010000010011010110010110111100101101100110100111101111101100001011110111100101010000; 
out4112 = 128'b00001100000010001000111100101011000000110010000000000101101101000011110110000001101000110100010000110111101110111001000111000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4112[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4112, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010001111000000110001001110101100011000100000011000000010000010000001010110001110001000000001010111101101111011011100111000; 
out4113 = 128'b11110111001010010001010100110000010000100000010010100110010110101011111100101011100000011011101001010110101011101010111001100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4113[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4113, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101110011000111111110111001100101000101111000000001110101010101011111010100001011111010111011100100000100001100010101111101001; 
out4114 = 128'b10101110110101100100001101101110100111010011101111000101101001001000011100000000000010011101100100111010010001010010110111100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4114[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4114, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011100110001111111101110011001010001011110000000011101010101010111110101000010111110101110111001000001000011000101011111010010; 
out4115 = 128'b01000010110010000100101101011001001011111110111000010011011000011000110011011011101001001010111011001100010000000101000110100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4115[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4115, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001100011111111011100110010100010111100000000111010101010101111101010000101111101011101110010000010000110001010111110100101; 
out4116 = 128'b11011101110101001110001001101001100000100100000101000000001110101001100110011111000101011011001010100111010110100010111111101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4116[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4116, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011000111111110111001100101000101111000000001110101010101011111010100001011111010111011100100000100001100010101111101001011; 
out4117 = 128'b11101111010010010100000001101100100100101011001101101011111111000100100001011010011100101001011001010010010000010010111011000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4117[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4117, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110001111111101110011001010001011110000000011101010101010111110101000010111110101110111001000001000011000101011111010010110; 
out4118 = 128'b00101101101001101110111010110010111100001010001111000010010010011001101111111000111111100001100100001111001011111000011010100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4118[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4118, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110011001000101110011000101100111111110000111101011111011010010101000100010101000101001001110011111001011000011100010110100; 
out4119 = 128'b10111110100101100011000000100000011110101100111000101000100101000001010001111111001110010010111111010100001000000101100001111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4119[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4119, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110110100110101110011011010111111100010001111101001011000001010101001001000010010010101000010110001101100010011010011110001; 
out4120 = 128'b11000111011011100100000001000101101010000000111010010010101110011111111010010111010101100100100011011101001100110011010001001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4120[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4120, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111101111010101110011100100001111011010011111101100011110111010101010011101100111101101011011101100100010110010110001111010; 
out4121 = 128'b00001010111001101001100100010011000111111011101000010110110001000011011100101101001101111101001110001110100010111010111001110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4121[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4121, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111011110101011100111001000011110110100111111011000111101110101010100111011001111011010110111011001000101100101100011110100; 
out4122 = 128'b11001111011110001011101101011110111001011011000110111111100010111100110101100000111010011011110000000110001100101011100010000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4122[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4122, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100111011101001011011000001001101110111111110001111010101000101010001111011011101110010110000111101110001011111010001110000; 
out4123 = 128'b10000111100001000011011000001100011011110100111010001011110100110101001010111000100101001011000111100011101100011011000000011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4123[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4123, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001110111010010110110000010011011101111111100011110101010001010100011110110111011100101100001111011100010111110100011100000; 
out4124 = 128'b00001011101111000110000010000010100100100000111000111100101011101111000110010110110001111111100100000110111010111011000101001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4124[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4124, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001101000011011111001010101000111000001111000000011111010111010111111100000110100001100011101111000111111101001010001011001; 
out4125 = 128'b01110001000000101100110101101001010010010010010001111011000111111000000001100001110101011111101011100001110101011001101011101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4125[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4125, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011010000110111110010101010001110000011110000000111110101110101111111000001101000011000111011110001111111010010100010110011; 
out4126 = 128'b11111100110011010111100101111010100110111001000101101111000000110111100101010100101100011011110100000111011110011010001110001111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4126[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4126, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110100001101111100101010100011100000111100000001111101011101011111110000011010000110001110111100011111110100101000101100110; 
out4127 = 128'b01100001010011101010110011110110111100111101011110110101001101111001000000100001011001000110100000101011010011000011011000111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4127[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4127, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101000011011111001010101000111000001111000000011111010111010111111100000110100001100011101111000111111101001010001011001100; 
out4128 = 128'b00111001101011111001101010010011101111101000110111101010110011000100111001001111111010011111011010010100010110001000001110100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4128[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4128, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101011011010100100000001110000111000010001010111110000110110111001100010111111110100001110110001100101100110101111011011100001; 
out4129 = 128'b01110011010010000010000001101100111100010011100011111000111001111010011110111011101101111011000110000000011001010110001000010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4129[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4129, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010110110101001000000011100001110000100010101111100001101101110011000101111111101000011101100011001011001101011110110111000010; 
out4130 = 128'b00111101011110011000010110100101000101011111001010001101001001110110000101101010111110001010000000100001010011001010110000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4130[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4130, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000110110000110100000110110011011001010100001000110011101101011111101001000000100100110101110111110011111100010010110101100100; 
out4131 = 128'b11000100000010110011010001011101010011100001011110101011100010111000001110010100001110111111110011110001011011011110101001010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4131[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4131, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100110111011001100001100010110001010111001000110010111101100000110110000111110111101100101011110000010011110001010110000101000; 
out4132 = 128'b00100011111010000100101001011110000000110111011000001111100011111100000001110101011011000110110010110111100011001111010000101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4132[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4132, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110101100111100011001011100101101100011011011011111101110110100000011000010001111000100001101100001011010111010111010110001; 
out4133 = 128'b10111010000000110111000000001011111111101010100010010100101101101101100111011000111011111100010011001000100111110011010110101110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4133[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4133, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101011001111000110010111001011011000110110110111111011101101000000110000100011110001000011011000010110101110101110101100011; 
out4134 = 128'b11111100100110010001001010010110100011111111000100111000111100010011000000000110110100010110101010101101101101101110100000011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4134[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4134, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001101001010101100100000010001110011100111010001110001101101001101110110111001000011110000111100000001101000100110000100110; 
out4135 = 128'b01101111100101001111000101100001100011111001001111011110001110110100101111101010101010011011001000010001111111100100001110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4135[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4135, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100011010010101011001000000100011100111001110100011100011011010011011101101110010000111100001111000000011010001001100001001101; 
out4136 = 128'b01101111010010000111000001111000111001010110101111010011100111100011110011110101010110010101001001100100011001001111000111100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4136[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4136, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101111111110010010001111000000001100010111111001000000000011111011001100011010101110110101111100101010010111100011001111010; 
out4137 = 128'b10000011100011011001000100011101011010110110111011110100000101100001111101000001111111111001111000001000101011100001011100101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4137[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4137, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011111111100100100011110000000011000101111110010000000000111110110011000110101011101101011111001010100101111000110011110100; 
out4138 = 128'b11101111101111100111111101001101001101001100101000110110111100110100101100101011011011011110000101110000001101010000101011101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4138[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4138, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111111111001001000111100000000110001011111100100000000001111101100110001101010111011010111110010101001011110001100111101001; 
out4139 = 128'b10010110100001110010101100101111011011011001011001001101011000011110011110111011101001110010010100110011100011100001011000100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4139[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4139, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000100100100110110001110110000110100000110101110110000110101000010101110100101011010111011001101001111110001001100010100110010; 
out4140 = 128'b00011011100010010001111010101110010011010111011111100110000111101100110110011101001000011011110000111110010110101100011011110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4140[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4140, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010010011001000011100010001010000011100001010010001011100111100111111110101000001111000101011111010000100110111110010000101; 
out4141 = 128'b01111101011111110110010010010100001111000011110011011110110010010111000010101000111100011100111100101010101100111110000010101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4141[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4141, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100100110010000111000100010100000111000010100100010111001111001111111101010000011110001010111110100001001101111100100001011; 
out4142 = 128'b01011101011101001011000111010001000101101001001111001111100101011110010000110101010111001000010011111011001011110010110101111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4142[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4142, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010010110000101110000110101111001100001111110110101000101001010011101101011110011101100011110001101110101110000010011110110; 
out4143 = 128'b01011000101111001100011001000010000100010000000001111100000100010001100011110010111110100001011100010111011010111011111011111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4143[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4143, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000100101100001011100001101011110011000011111101101010001010010100111011010111100111011000111100011011101011100000100111101100; 
out4144 = 128'b01011110110111010001000100110100010001011010000010101101110000100001110001011001100001000101001111011111110111001101101101100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4144[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4144, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010000010110011000010100111011110010110101100100100100010010000010100010000111010111111001001010010110001101110010100111000; 
out4145 = 128'b00100111010110010001101010101110000010110110100100111101010110100010111001101101011011101101111000110010001101000111011100000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4145[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4145, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111011111000010000100111110000100111100001110111001110010011001001010011110000001110000100011000000000101110011110010010001; 
out4146 = 128'b00000100101001100101110000111110000001001010010011110011001101010110111111101111001110000100000111110110110010101100111011000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4146[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4146, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110111110000100001001111100001001111000011101110011100100110010010100111100000011100001000110000000001011100111100100100010; 
out4147 = 128'b10100110101001111001001111010000010101111010101111000010001111010100100110001000100110000101110011101110110110001000111100111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4147[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4147, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111101111100001000010011111000010011110000111011100111001001100100101001111000000111000010001100000000010111001111001001000100; 
out4148 = 128'b00001111011111010011010101100010001100001011111111101001111001011100100000001111100001001000000100001000000001000110100010100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4148[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4148, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011111000010000100111110000100111100001110111001110010011001001010011110000001110000100011000000000101110011110010010001000; 
out4149 = 128'b01110101111110010011001100001101110110111110100001101000010111011100010010101111101011100100100100101001100001000001010010010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4149[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4149, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110111110000100001001111100001001111000011101110011100100110010010100111100000011100001000110000000001011100111100100100010000; 
out4150 = 128'b01111101110110100010010011001101111010011000111000110100001100100100001101011101101100001100001010110011110001011100111111000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4150[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4150, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000100111011100110011110110010100110010110001011001001111010011100101101111111001100011111010001100111011111010110010011000000; 
out4151 = 128'b10100111111011111110000100010001101011111010010011011100011100011001001101000101111111001000000110011101110011001001111010101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4151[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4151, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100010101101101000111100010101110100111101000001100011000010000000111001000001101100110000010010101011011000000011111101100000; 
out4152 = 128'b01110100110111101111001001100011100111010010101101110010111001100010101010101111001001101000100001001000000001100001100000111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4152[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4152, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101110000001110101111001011011010001101011010100110110110010111000010000111100101101101110010100110011010110101000100000100000; 
out4153 = 128'b01110111001001110011011001110110010111100111110010000001010000001000010111100111010000100001001011000001111000010001110111011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4153[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4153, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100000011101011110010110110100011010110101001101101100101110000100001111001011011011100101001100110101101010001000001000001; 
out4154 = 128'b10111111110000010110001100000011011010010001010100100001010100110101010110111100000001110110011000010111000000001101011111111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4154[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4154, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010011011101110011100100011101111110111100000100101011111101011000100001001101000010110111100010101000111100001101011001100011; 
out4155 = 128'b11110001010010010110011100011011010010010011000101000111010001101101110001011110101101000101011010111011010011001000000111011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4155[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4155, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100110111011100111001000111011111101111000001001010111111010110001000010011010000101101111000101010001111000011010110011000111; 
out4156 = 128'b01000101011000000011010100011100100000110000100110100110000001110110011101001011011111111011011111111011111101011110101100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4156[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4156, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100110101101101010010000000111000011100001000101011111000011011011100110001011111111010000111011000110010110011010111101101110; 
out4157 = 128'b00100101101110100111001011111011010111000001110001011010001010111110011111110101011001110010000110000100010000001001101110101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4157[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4157, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001101011011010100100000001110000111000010001010111110000110110111001100010111111110100001110110001100101100110101111011011100; 
out4158 = 128'b00110110001001100100011110100111100100100001110100100111000110010111110010101011011111011011110100010011010110001010101110001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4158[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4158, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010110110101001000000011100001110000100010101111100001101101110011000101111111101000011101100011001011001101011110110111000; 
out4159 = 128'b00100101110101000011000011010001010100101011100110011000001000101000111001111010101100111001001101011110000011110100110011000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4159[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4159, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101101101010010000000111000011100001000101011111000011011011100110001011111111010000111011000110010110011010111101101110000; 
out4160 = 128'b01011000001101101010010101011011001011011110010101111100110011110001011111100000011011100001111011101100001010110000111101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4160[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4160, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110000101111110011001001000000011100110100010000001011000000110010101000001110000101001000000101011011111101111111011000011; 
out4161 = 128'b11000001010101001011100011011011101111001001101001110111111111110110000101101101010010111110011000101001001001000011111100110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4161[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4161, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001100001011111100110010010000000111001101000100000010110000001100101010000011100001010010000001010110111111011111110110000110; 
out4162 = 128'b01111100011000101111100100110110111110011110011000110110010100110001000100001111011100011010111010101000011111100111010000001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4162[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4162, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110010010000111111101101000001101111100101010000100111000011111000001000110110010001101000010000110100001010000010111001111; 
out4163 = 128'b00010111011101001110100100001100101001100011001100010110111011011000010011111001111000100100101100000111001001110000011100111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4163[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4163, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111010100001110001100010011000011000011111110110001000101000111000010111001100010100110011000100100110011101001111010101011100; 
out4164 = 128'b01001101011110111111011010011001000100110110000111100001001001101011011011000001011100110110001110101010010111100001110110100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4164[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4164, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011000110011101011101111000110011011001001110010000001001110110111011011001011001001111001001100111100101110001010001111011; 
out4165 = 128'b01001010011100111000010000010001100000001010110111110010110101110100110111001010001011101100001011110111011111111001001001111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4165[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4165, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110001100111010111011110001100110110010011100100000010011101101110110110010110010011110010011001111001011100010100011110111; 
out4166 = 128'b10010010111001110000101101001001010010001100101000000011001001010000111011000111110101011111001000100011110110100110101001110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4166[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4166, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001010011100001011101110101011001110000010011011000001111111011101111000100100010100010101100110110101001000101010111100101101; 
out4167 = 128'b01011110111010001010100110000100101100100100110111100111001011111100111101111100011001100000010001110010001000110000110010000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4167[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4167, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100111000010111011101010110011100000100110110000011111110111011110001001000101000101011001101101010010001010101111001011011; 
out4168 = 128'b01011111010101010111000100000111011110111110011001100011010000111101101110010001100011101010010101101001000000001110100100101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4168[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4168, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101111110101010000100011100100111011101111001110000110100101110001110111010000100001111111011011111111111101000100001001110101; 
out4169 = 128'b11110110110100010000001110100110001011101011111110110111010100110110111100101101100100000001011110101011001101011011101001010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4169[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4169, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011111101010100001000111001001110111011110011100001101001011100011101110100001000011111110110111111111111010001000010011101010; 
out4170 = 128'b10111101001001000100111110111001011101110111110011101010010100110010011101000111100110100111001110101111111101101010011101011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4170[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4170, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111111010101000010001110010011101110111100111000011010010111000111011101000010000111111101101111111111110100010000100111010100; 
out4171 = 128'b10110100100101101000000010010001101101110001101011110101100101000010011010111100111110000100011000000000011001011011001101010101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4171[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4171, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111000101111111010000101101111011110011111010010110101110110001000101111000101111111010010011111010100110111001110110101101010; 
out4172 = 128'b01000010100110101100001010001010110111010101010011010101100100001100010000110010000111110111011000101110111101011100000100011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4172[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4172, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111011010001010010010010110111111011000000111101010110100010111001011001010001110001101111110000010110001110010010000010111; 
out4173 = 128'b10110100111110111010010110010101001101010101100100001110111100010111101110110111110111110000001101000011111111001010101000100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4173[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4173, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101110110100010100100100101101111110110000001111010101101000101110010110010100011100011011111100000101100011100100100000101111; 
out4174 = 128'b10100011000000011000111110010110101001100000100100000000110010010110001111000010001100101000110011100101111100001100001000100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4174[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4174, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011011101101010111010000010011111110000110111100101010001001011010111001101001001000011110111000100000011000100110111010011101; 
out4175 = 128'b01000111001000001001100000111101100111001010101101101111101101001100100101100100011010001001000011100100110110111100010101111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4175[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4175, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111011010101110100000100111111100001101111001010100010010110101110011010010010000111101110001000000110001001101110100111010; 
out4176 = 128'b11101111110010001001011101010010110000011001010010100000100001001000101101100010001000111101100010010010110001101001001100110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4176[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4176, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000110000100011011000000111111011111101010000101001111101101101110011100101010001010010100010101010111101110100010010110111; 
out4177 = 128'b00001011010111101111110001101100000111001111001110100100000110000110110111001100110101101001111011001101001001110001110101010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4177[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4177, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111100100111000101001000111110100011100000011010010100011011101110010001011010010001100000101111110100100000111011110101101; 
out4178 = 128'b11010101110110000010000111100010101001011101011011010001101001011101001000101001110110110000011000000110111011000100000101000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4178[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4178, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101111001001110001010010001111101000111000000110100101000110111011100100010110100100011000001011111101001000001110111101011011; 
out4179 = 128'b00100111000111011111010110001111001101000011010011010010010011001111101101010110101110001011011001011111001111011010010011111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4179[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4179, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011110010011100010100100011111010001110000001101001010001101110111001000101101001000110000010111111010010000011101111010110111; 
out4180 = 128'b10000011001010000011110110011110001001011010010010010100110000001100100001000000111011011111011111100101110001000100001111110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4180[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4180, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111100100111000101001000111110100011100000011010010100011011101110010001011010010001100000101111110100100000111011110101101110; 
out4181 = 128'b10111101110101010100010000111001000001010100011111000101001010101010100001101001110001101011001101010100001001001000100011011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4181[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4181, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001001110001010010001111101000111000000110100101000110111011100100010110100100011000001011111101001000001110111101011011101; 
out4182 = 128'b01111101101010100001110001101101010010111110101100000001101110010000101111101011000100000111110010000000000111010111011101000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4182[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4182, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110100011001101010111010110010001101100111001011010000110110111111010000101000110110101011111111111001011100000000101101111001; 
out4183 = 128'b00000001011110000011110111011110100101101110111000011000100100100010011011010011100101000101000001011001111110100110011010000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4183[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4183, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101110110110101011101100101100011000101000110100100000110101111000110100010000011101111110111111011001100111101110100000110000; 
out4184 = 128'b11010001101001111000100010100100101011010100101010010000000110110110011000001010001001010001100000001100101010100111100110011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4184[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4184, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011101000101001000000010000110010110111001011000000110011110111111101100001001011010100111110011000010000110010111010100010; 
out4185 = 128'b00000010000010101100000011001011001010001000110111101000101110110011111010100010100101011100110000100011100100101111111101010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4185[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4185, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111010001010010000000100001100101101110010110000001100111101111111011000010010110101001111100110000100001100101110101000100; 
out4186 = 128'b11000100011101100000011001101000101010000011010001101101101010100101010101011101001101011001000110100011011110001000000011010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4186[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4186, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101000100111011010011000001011001000111010001110000010010111011001100011000101011101111010111001001010011100100100010001001011; 
out4187 = 128'b00101010111110101000010010011000010101110011111101010010000100010100011001001001011001000111011110101011101110100001001111000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4187[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4187, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010001001110110100110000010110010001110100011100000100101110110011000110001010111011110101110010010100111001001000100010010111; 
out4188 = 128'b11101000101001011010000100001101011000100001000110010101100010011101010111101111001110101101110100100001100110011000100010110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4188[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4188, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100011000010111111001100100100000001110011010001000000101100000011001010100000111000010100100000010101101111110111111101100; 
out4189 = 128'b01101011010101101011001111000101001011111111101110110010000110110110001100000011111010001101110100011010011110011011110000010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4189[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4189, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001000110000101111110011001001000000011100110100010000001011000000110010101000001110000101001000000101011011111101111111011000; 
out4190 = 128'b11101000010010101010010101001101001000010100101010001010101110101101101001100010110111100100000010011101011110101111001010010100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4190[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4190, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010001100001011111100110010010000000111001101000100000010110000001100101010000011100001010010000001010110111111011111110110000; 
out4191 = 128'b00010010010001000010001011010111011001110001000011101101110110000111101110010010111111001101010100000110101111000000110100111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4191[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4191, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100011000010111111001100100100000001110011010001000000101100000011001010100000111000010100100000010101101111110111111101100001; 
out4192 = 128'b00100100110000111000001001110010101101001010101100110101100010011011001001111101010110001101100010010110010100011110001100001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4192[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4192, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110110011100011010110000100100011101000101010101101011001111100101010110111111110110010011100011000101000010101001001111100111; 
out4193 = 128'b10100111110001100010000111001010001110110101000000110100100111111000110110101100111011111101111011010000011110001001010110100001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4193[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4193, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100111000110101100001001000111010001010101011010110011111001010101101111111101100100111000110001010000101010010011111001110; 
out4194 = 128'b00110100111010011111010001011110011101101110011101000000000001100100111001011111100101001001100101110110111010100111011001001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4194[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4194, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111101101110001110010110101101001010000000011000111110001110000001101000000101111011101101111010001001000001101110001111011; 
out4195 = 128'b10110111110111011100010111101011010010010110010010010100111000100111010111110011111000011010101110110110111010000110100100000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4195[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4195, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001000111111001010101001111001111100101010011100100101100000101001100111110101000101000111101100111010010110010101100010001; 
out4196 = 128'b00110001010010101011110111111110111011101101010000010111100111111110101100110010101110111010000100111000101001101000111001110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4196[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4196, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100100010011101000011010111010000010001111110010100010010111101111001111000010100111000010011000001011100111001100010111000100; 
out4197 = 128'b11010110110001011101110110111111100011101101010010011011100111110100110011010000101001000100001000111111100010111111010000111011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4197[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4197, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001000100111010000110101110100000100011111100101000100101111011110011110000101001110000100110000010111001110011000101110001001; 
out4198 = 128'b00111001100111100110110111101100100110111010011100011110110111100110110010100000101110110111001111101100111011011011011000001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4198[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4198, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111010010111011011011001100010101111010011111100010010001011001101010110101101010011010000011101011011110011000010011110100; 
out4199 = 128'b00001110101011111010010011111111001000001111110010011101110111100101111110101110110000011110001001100111001110101100101010101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4199[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4199, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001110100101110110110110011000101011110100111111000100100010110011010101101011010100110100000111010110111100110000100111101001; 
out4200 = 128'b00100010000101011111011111000010010001001101010010101000110110011001011111010010110100000010110010001110101100001111101100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4200[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4200, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011010111110111011100010101001010101100101011100010001010000011111101101001011111111011101101101000111011001000000000110101; 
out4201 = 128'b10110001111110010001101101001011000010011011010010000100110011110110000110010000010111101001000110110101110100000010010100001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4201[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4201, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010110101111101110111000101010010101011001010111000100010100000111111011010010111111110111011011010001110110010000000001101011; 
out4202 = 128'b11011001100011110011011011111000101100111110000101000101011100110100000111110001000011010000001101101111110111001111100110100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4202[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4202, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101011111011101110001010100101010110010101110001000101000001111110110100101111111101110110110100011101100100000000011010111; 
out4203 = 128'b01101111010011011001101001100110110000110011000010001111001110110101100010110110011001101011101111011100001010011100001110010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4203[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4203, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101100100010100001010010001101001000100000001001111010011111111010111011110100001001001110001110000010011011101001001001001000; 
out4204 = 128'b11000101001010101010001101001000110111001101101110110101101010111010010010101000001001011000011101011101001110101011100000000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4204[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4204, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101111011001011000010100111110001100000101000110011111110000010000100001010111100100001111111111000001110101111011011101110111; 
out4205 = 128'b10011000010011101101100010010111110010111100011101111111011100100100101001101010010000000111101001011000110011010001000000111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4205[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4205, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011110110010110000101001111100011000001010001100111111100000100001000010101111001000011111111110000011101011110110111011101110; 
out4206 = 128'b10110100010101100010011010101100011101011110110011000011011011000001100110011110000011001101110011011110111011111100001110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4206[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4206, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011111001111011100011011100101101010001001100010100001110100111010011100001100110101100011111000010010101000100111000111010; 
out4207 = 128'b01011010001011110110000011101011010110101101101011010100111011111000100000110111011101010110100100001101111100111111111110100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4207[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4207, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111110011110111000110111001011010100010011000101000011101001110100111000011001101011000111110000100101010001001110001110100; 
out4208 = 128'b11100101100101010110101010101110011111110000000100000010110000011011111111101110101011010011111100011101010100001101011010101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4208[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4208, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011001111011110100111101010110101000000001100100111011110101111000011000111001101100100010011111001100010110111010101100001111; 
out4209 = 128'b00111000010001111110100100101001100111011010000001100111101010000011011000110110000011100101101100110110000101001111100110100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4209[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4209, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101101011110011001010001001001101000110011100011100100100010101100111001100101111010111011101011101101111011100010111111001; 
out4210 = 128'b10111110100110001001000101111010100010010001100111010101000100010100100001111010010000100010010111001110101000010110010101100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4210[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4210, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011010111100110010100010010011010001100111000111001001000101011001110011001011110101110111010111011011110111000101111110011; 
out4211 = 128'b10000100100111100101111000010101001000010001000001111000011001010000011100000001101011001001111110111010111011010101011100101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4211[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4211, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110101111001100101000100100110100011001110001110010010001010110011100110010111101011101110101110110111101110001011111100111; 
out4212 = 128'b11100110100100000000000001001010000000111101110111011110011001110001001101001111110110111010111011000000101101111010000000100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4212[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4212, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101101011110011001010001001001101000110011100011100100100010101100111001100101111010111011101011101101111011100010111111001110; 
out4213 = 128'b01001100110010001101010101111111101001011001110010001110011110111100001101010010001110000010111111000011010111010011110100011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4213[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4213, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011010111100110010100010010011010001100111000111001001000101011001110011001011110101110111010111011011110111000101111110011100; 
out4214 = 128'b11100100110111110100110010011000001110101010000000100011101010000111001101101111010011110010011101010000001000111101100001000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4214[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4214, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000011100101111111110100000010111110001011011011111001000101010110110000101000011101111101001101110010101100100010110011011111; 
out4215 = 128'b10110011111000111011100111110110000001101110101110111101101100101101100010000001001111110011011111100000000101000101101001000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4215[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4215, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110001010111100101011000100001100001010011100010011001000101001000110111101111001101101001111000100000011011101100101001011001; 
out4216 = 128'b00001111011000000010111101111000001111010000101000111001101000011110100101100010011110110000111000011011101011101100111100110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4216[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4216, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100110011010000000001100111011111100010010001011001000101110100111001100001101101000000010010000101110101110000011101010100; 
out4217 = 128'b11100001000011011001100001111101001011010110011000000101001100000011011011101010111011111010011010101101011000010000110011110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4217[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4217, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001100110100000000011001110111111000100100010110010001011101001110011000011011010000000100100001011101011100000111010101000; 
out4218 = 128'b10000110001010111100111100100001010001010101000110011100100000100000000010111110000111011011110100101011101001010100101000110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4218[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4218, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101010001011010110110111001100011001100010000001111011000110110110000111001000010010010101011010010010101101000111010110110; 
out4219 = 128'b10110010101001001100100011101001011110110000100100011000110010001101010101110000010000111001110001011111101000000101001000101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4219[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4219, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010100010110101101101110011000110011000100000011110110001101101100001110010000100100101010110100100101011010001110101101100; 
out4220 = 128'b11001110100101010101011011000000101111001110110000101000000110100101111111000110110101011111000011100110011111011110001011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4220[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4220, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100011011001110001101011000010010001110100010101010110101100111110010101011011111111011001001110001100010100001010100100111110; 
out4221 = 128'b01100010100110011000100010101110111000010111000100110101100011111000010111100000100001111001111010011000001111000010011000100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4221[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4221, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000110110011100011010110000100100011101000101010101101011001111100101010110111111110110010011100011000101000010101001001111100; 
out4222 = 128'b00110101000101101100101110000000101100100111000011100000101000011111011111101001101110011001100111011010001101001110101101100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4222[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4222, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101100111000110101100001001000111010001010101011010110011111001010101101111111101100100111000110001010000101010010011111001; 
out4223 = 128'b11101111100111101010100011001001101000111001011010101000000111100110110001100111001100001001010010011000001000101111110001011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4223[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4223, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011001110001101011000010010001110100010101010110101100111110010101011011111111011001001110001100010100001010100100111110011; 
out4224 = 128'b11111100100100000010001100110001101000101111010001100100101011110110011011110011010001000100010000100110111111001111010111101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4224[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4224, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010101101110010001001100001100011001100011001111101000101111101111101101011000011010010010001000010011010101110000110010001011; 
out4225 = 128'b10101111010101100010010011101100011000010001101111000000010100001101011011001100001100110011000010100000101010010010000100111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4225[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4225, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101011011100100010011000011000110011000110011111010001011111011111011010110000110100100100010000100110101011100001100100010110; 
out4226 = 128'b11101010010100111001110111000011000110001110101111011001010001010100110100111100010011011001011100010110000110010000101010011001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4226[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4226, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000011010111010101111100111101111111101111110001001010010001010001011000111001110011011010101001011110000010110011111010100111; 
out4227 = 128'b10011001110010011111110101000111010001000110110111001111011101101000110011011001000111101000111101110111111100110101100110011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4227[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4227, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010011000000111010110101110111100110111100101101111100001101001101011100101011111100100111011010101111010000010111000111000101; 
out4228 = 128'b00001011000100010000111000101101101110001101011001111011011011001110000101000001011011101110100110111110000100010011000001010111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4228[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4228, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110011101111100100100111100011010100011010010100010000110101110101010100001111100011011100111101001101110101011110111100000001; 
out4229 = 128'b01010000011000101110100000000100101010011011100010101101111101110010111101111110001101101100011111100011000000111110000100101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4229[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4229, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100111011111001001001111000110101000110100101000100001101011101010101000011111000110111001111010011011101010111101111000000010; 
out4230 = 128'b11101010111001010101001000100101101010101001001000101010100010000101010000100001011011000000100000100110101110111001010010111110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4230[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4230, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011011010000000011010010000001001000001010011110101011111000111010111101100110010111100001111100100100000000001011000010001111; 
out4231 = 128'b10110101111111101111010110100101010110101100001001111101011001010111101001111001001010010001100011111111010011001100011011000101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4231[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4231, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110110100000000110100100000010010000010100111101010111110001110101111011001100101111000011111001001000000000010110000100011110; 
out4232 = 128'b10111010001001011011111111110010101011010010111101100011110000000101110100111001111100011011001101011010011000101010011101111000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4232[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4232, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111000101110011100000100001000111001001010110101000111001100000100011011000001000100010101111010000011010101011100111010110111; 
out4233 = 128'b10100111011001000011001111110111111100000111000001011010100111001010000011110011101001001010111000110111110001011010111101111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4233[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4233, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110001011100111000001000010001110010010101101010001110011000001000110110000010001000101011110100000110101010111001110101101111; 
out4234 = 128'b10100101000001000101011011100110010000000001100100100000100011010011100010101001001011100110100010011101110010001111100110100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4234[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4234, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100010111001110000010000100011100100101011010100011100110000010001101100000100010001010111101000001101010101110011101011011111; 
out4235 = 128'b00101100000011111011100000100011010000111110010011110101000001001000111110110000110100100010001110001101000010000110011110011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4235[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4235, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010000011101110001101101001011010000110101100111010001001111001100110101010000111000111101011000001001111110010111100100110100; 
out4236 = 128'b10011000010010000000011011001111001100100110010001001000100011010100000101100011110100100011001101100110010100001010110100100100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4236[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4236, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101010101110010010110011010111000001000000001001010110001110110000111111001101011101000111000000000101001011111111011100010; 
out4237 = 128'b11100110100001101100110000010100000110100111011011110011111010101100111111010000101101011011101100010000111100010100100101100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4237[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4237, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010101011100100101100110101110000010000000010010101100011101100001111110011010111010001110000000001010010111111110111000100; 
out4238 = 128'b10011110011001001100110000101110101000011111111000100110001001110010111001110010100001100011011110100111111001101100000100010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4238[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4238, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000000111001011000010101100111111001000011001011000011101000110111110010111110110100110001101000010001110000001111011100000011; 
out4239 = 128'b10100001111011011111001001100100001011000100011101000000000111110110001010110011100110111011101001111001011001110111101001110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4239[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4239, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001110010110000101011001111110010000110010110000111010001101111100101111101101001100011010000100011100000011110111000000110; 
out4240 = 128'b01101110111011101111110001000010110111011011001001010111001110010110001010011110001100100101111110010010011001001110001110110110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4240[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4240, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10010110001011110000011010010011111101101111100011100110001100110000100110100011001001010100101001010100010101001101000010000110; 
out4241 = 128'b10100111100011100001010101110101010000100000000000100001101001100101011011111011100101101011101011001001111100010100011011000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4241[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4241, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001111001110001111000101011100010111100001000100100110110001110100000011110001000111011011010111011111111101010110110000110; 
out4242 = 128'b01000011001110110010001010111000100111000001001011110000011001110000100011110011100001011100100100111101010110010110010101100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4242[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4242, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110011110011100011110001010111000101111000010001001001101100011101000000111100010001110110110101110111111111010101101100001101; 
out4243 = 128'b00000100011001111110110110101111011010111001000101100111011011100111100010110010000111010000010111110111001100101110110101001010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4243[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4243, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100111100111000111100010101110001011110000100010010011011000111010000001111000100011101101101011101111111110101011011000011010; 
out4244 = 128'b11010001101110011100010101110101001100010011001010101100010010001001100010000100011000001011010010100110011110110010000111000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4244[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4244, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001111001110001111000101011100010111100001000100100110110001110100000011110001000111011011010111011111111101010110110000110101; 
out4245 = 128'b10110010010110111010001111000000111111010110010111010110101000110011010110000001101001010100011110110010001011100111110100011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4245[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4245, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011110011100011110001010111000101111000010001001001101100011101000000111100010001110110110101110111111111010101101100001101010; 
out4246 = 128'b01000111110011100011101100010111111110001001111110011100001011010011000111011001000100000100111110111111000000110111001011100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4246[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4246, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101001010110101101011001111101000111100111011101110011101000111111100010011100000111111111010101101100100000101011110001011110; 
out4247 = 128'b10011110111010111011010101100010001001111010000111110101001011011000110100011101011011000101001000101100010010110010111110000110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4247[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4247, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000111000011001011111111110110010110101101110100001111111110010000101001100000010101101100100011001010010100100111010000110110; 
out4248 = 128'b10101000011111100100111100101111011001101001111000111000001110010100010000110011111011001101001001000110010010010111111010011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4248[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4248, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00011011101000000110110011100000110100111000100111110111010011001110111110011000110001001011001110000111111100111110010011100110; 
out4249 = 128'b11010010010101110001010001110001110101000011111011010000111110111010111001010101001001110101111101111100100110011000010001011000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4249[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4249, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110111010000001101100111000001101001110001001111101110100110011101111100110001100010010110011100001111111001111100100111001101; 
out4250 = 128'b01111101110011010011001001100001011101011110000000111001110000001000101101011101011010000110101000011001101100010000010011110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4250[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4250, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011001110001010000010001111001010000001010000110101100011010100010100111011011110111110110000001100100110001001111100010000; 
out4251 = 128'b10000000110101000110110000010110001111110100011000111110110110010111010001000100000100011001000110110011100010010001001010000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4251[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4251, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110011100010100000100011110010100000010100001101011000110101000101001110110111101111101100000011001001100010011111000100001; 
out4252 = 128'b11111011000011111000101011111000110100100010011000111111000011011110100100100111011110000111000000011011110111110010011101000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4252[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4252, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111001010110111001000100110000110001100110001100111110100010111110111110110101100001101001001000100001001101010111000011001000; 
out4253 = 128'b10000111011111111100000100101111010011000001001111000011010110100111111000010011100011110011010111000000011101100000101010000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4253[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4253, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110010101101110010001001100001100011001100011001111101000101111101111101101011000011010010010001000010011010101110000110010001; 
out4254 = 128'b11110111100010101110001011111110101111001001010111001011000100000010011011100000111101100101000001110011010001110000001110101100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4254[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4254, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11100101011011100100010011000011000110011000110011111010001011111011111011010110000110100100100010000100110101011100001100100010; 
out4255 = 128'b11010001110100111101000110001010100101110001110001001011010010101111110001110111110000010001100100101111011000011111111101011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4255[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4255, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001010110111001000100110000110001100110001100111110100010111110111110110101100001101001001000100001001101010111000011001000101; 
out4256 = 128'b11000110100101011101101101101110000101011011011110000100000111010000010101101111001011000000000010000010110100011111100001001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4256[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4256, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101111101100100010010000010011000011100110011001000001101010011101011010110111101111001111111001100010010101100010001001110010; 
out4257 = 128'b10010101001110000111110000000111110011100110000101101111000101110001101110000110100110011001000010001010101110100110001001110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4257[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4257, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011111011001000100100000100110000111001100110010000011010100111010110101101111011110011111110011000100101011000100010011100101; 
out4258 = 128'b10010100110100011000101101011001001001010100111011010101111010101000110110011100100001110010111111000011111101011100000001000010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4258[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4258, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001011110101011010001011111001101111111111101000111000011101000110001101001010011110000011111101011000011101010101110111001; 
out4259 = 128'b10011111101011001110001110110011000100000010101111010100110110011111111100101010111100011110000111010111000001001100100010001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4259[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4259, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001101010001110100110010101101011000011001100011001111101101001100111001100101001000101111000110110100010010110111010100000001; 
out4260 = 128'b11001011100001110011110111111100100000010111001001010110010111011101010111000000000101101011010100110111100111001001110010101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4260[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4260, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110101001111001011110101001001110011010101011111011110110000000100101001111101111110010001110100001010110000001100100001110001; 
out4261 = 128'b00101001011011100011101100011010110011000101100110011101010111001001111010010010001110001010100100110000101001011100001010001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4261[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4261, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010011110010111101010010011100110101010111110111101100000001001010011111011111100100011101000010101100000011001000011100011; 
out4262 = 128'b01101111101010001100011011101110001010110111101110100000001111100010101001101100000110100010100000101001111001100001010000111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4262[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4262, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111011010000001101000100110100001110110011100100111010101010001111111101000000010110001000101001001001010101010000001110110100; 
out4263 = 128'b11101011100011110101001100000001001011110001101111100010000010010111000010100110010001100000010001001101100101011010111001101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4263[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4263, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110100000011010001001101000011101100111001001110101010100011111111010000000101100010001010010010010101010100000011101101000; 
out4264 = 128'b01011000011100011100111111101110000000011101001010011101111100101110001010110110001001110111100010000110000111111111101110011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4264[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4264, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000010101100010110000011000011111000101000001010101011000010100010101110110110110111101101011101000111000000100010110010100011; 
out4265 = 128'b10110100011111100100010100010101111101111101111010100101001010101000110000100100111110110000011110001001110001000011101110110111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4265[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4265, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000101011000101100000110000111110001010000010101010110000101000101011101101101101111011010111010001110000001000101100101000111; 
out4266 = 128'b10101000100001110011100101111000111011111101000000111101111000101010110100010111011001010010101000000100000011101000111011010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4266[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4266, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001010110001011000001100001111100010100000101010101100001010001010111011011011011110110101110100011100000010001011001010001110; 
out4267 = 128'b00011101110010001000011101110110110000010111000110010010111010100011001111000010011100100011010010100110000101001101101110101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4267[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4267, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111010001110010010001000001100000110100111001100011001111110001000101100000001010010100100010001011010010001110100011101101111; 
out4268 = 128'b11010001011010010001110101001010101101000010100010100101000000011001100000001100110001100001110101110001010100011010111110110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4268[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4268, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11011011110000000110000000001011001110101000000001110010010110001100000010110101001010000111011011010110110110001010110010101101; 
out4269 = 128'b10010011100011000010101001001000010010001110101000001010001001111100011110101001101101101111010111100110001110100010001011001000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4269[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4269, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110111100000001100000000010110011101010000000011100100101100011000000101101010010100001110110110101101101100010101100101011010; 
out4270 = 128'b10110010010010110110000000011100011000011110101010010111111100101000110111111010000000100010000110001001001011010011101111000001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4270[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4270, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000000101100111010010000111111111001000110011110001000110010101101010001100011000111010010010100111001001101001001000011000110; 
out4271 = 128'b00001000000110100011010111110010011010110000000000001011010001110001010111100001001111001111111110110011010100000110101001110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4271[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4271, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000001011001110100100001111111110010001100111100010001100101011010100011000110001110100100101001110010011010010010000110001100; 
out4272 = 128'b01101110001001111000011101000010010000010000010001111001010000010000011100100011001110001001000100111110001101100100011011001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4272[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4272, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101101011111001011010011101100100111111111100001100010100000101000011100111011110010000110101010000110100001000110000101101010; 
out4273 = 128'b01110000011000001000010000100110010101101001110110001100101100001111010111010011100100110010010001111100101011110110100001000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4273[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4273, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110101010010110100110111001010001100011001011010000100101011001101100011000000001011000010101101101111010111101110000010100111; 
out4274 = 128'b10110000001111101110000011101110001111001111100011101100100111011000000000101011011001111100011011101010110100101010111100011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4274[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4274, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101010100101101001101110010100011000110010110100001001010110011011000110000000010110000101011011011110101111011100000101001111; 
out4275 = 128'b00111100011001010000110111001010111000011110101000010001010110100111001110110111111011110001010111011110110111111010010000010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4275[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4275, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101001011010011011100101000110001100101101000010010101100110110001100000000101100001010110110111101011110111000001010011110; 
out4276 = 128'b01110000111110001101001100001101111000010001001100010000011101101101010101110010110011100101101101110010110010011111100111010000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4276[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4276, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010010110100110111001010001100011001011010000100101011001101100011000000001011000010101101101111010111101110000010100111100; 
out4277 = 128'b01010101000110010000111011000101001011100111011010001010110011011001101110011100100010110110101101011001111101000100010110001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4277[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4277, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100101101001101110010100011000110010110100001001010110011011000110000000010110000101011011011110101111011100000101001111000; 
out4278 = 128'b11101001101111011000000111011111001011001101100010001101001100110000100110000011001000000001001001101110011000100111000001110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4278[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4278, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000110110110111001110101010101001111001011011011010100001100101100111010110010001110011001001110001001100010100011011010000011; 
out4279 = 128'b00001111001011110101110101101111011000011100111010110001000011011001010111000100001000001011111100001000100001101000011110100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4279[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4279, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100010000001010001111010111001011101110000101111101001110011000100101111010011110011111101100101110001010000100100111101110101; 
out4280 = 128'b01010111001000100100110000110011010101110101110101011111101100000011000000000000111110101011100001001010100101111010110001001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4280[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4280, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101011101110000001100101100001111000000111000110010010001100010100000100010000001000110100110010000000110100101011110010011001; 
out4281 = 128'b10010111000101010010000000000110000000100011110110110001101111111101101000111111011111011001110111011001000000111000100010011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4281[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4281, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010111011100000011001011000011110000001110001100100100011000101000001000100000010001101001100100000001101001010111100100110011; 
out4282 = 128'b00011011100010010000001001011001010101000010000110000101011000011101010110110110000101100000000010001011111001011100101100101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4282[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4282, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001010100100100000110010100100011111010000000001001011011001101001011110111001100011100110001100001000111001101000000010101; 
out4283 = 128'b00110001011101101100101110011000000101110010000100001001011100111011010100000110100011110011001111010101110111100100101001110001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4283[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4283, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010101001001000001100101001000111110100000000010010110110011010010111101110011000111001100011000010001110011010000000101010; 
out4284 = 128'b00110011010111111111110000100010001110101110100001101110011000111111001111010000111110011111010110101101010100111000101001011111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4284[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4284, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101010111110110010001001000001001100001110011001100100000110101001110101101011011110111100111111100110001001010110001000100111; 
out4285 = 128'b11010011011110011000100101101010101011101111111000111000111100111000110101111111110101110000010000011111100010010111001011101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4285[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4285, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010101111101100100010010000010011000011100110011001000001101010011101011010110111101111001111111001100010010101100010001001110; 
out4286 = 128'b00011110100010101101000011101101001110111011000001110101100100101001001101001010110111100110100000101100111000111110010001010010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4286[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4286, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10101011111011001000100100000100110000111001100110010000011010100111010110101101111011110011111110011000100101011000100010011100; 
out4287 = 128'b00001001101001001010110110100011000111100000001000000101100101101110100011001110000010001111100101001101110101001101001000111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4287[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4287, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010111110110010001001000001001100001110011001100100000110101001110101101011011110111100111111100110001001010110001000100111001; 
out4288 = 128'b10100010100111010110101110010100010000111100101010011011100010010100111000100010000101000001101100010010000110110101100110011110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4288[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4288, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01101010110000011101010011011000100010011010000110001100110010000100011101100100111100101110110011011010011100101011110110100000; 
out4289 = 128'b11111000011110110011100110110010110110010111101000001011000111001001001000111000111100111100010100101011000111010110101101111100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4289[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4289, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11010101100000111010100110110001000100110100001100011001100100001000111011001001111001011101100110110100111001010111101101000001; 
out4290 = 128'b00110100101110101001010110001101100011111010001000001100100111000001001110101001010101101111110110010100100100001111110010101111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4290[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4290, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000001110001101000011110111010101011110010011110111111111010010101101011110111001110010101111110110011101110000100101100100011; 
out4291 = 128'b00110011010111001010010000010001001011011111001011011111001110001101011110001101111001111100000000111001000111010011000101011011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4291[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4291, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001010011001101101110101101110101111110111011110011000110101111001010001010100000000101001110111101000000100010101111100111; 
out4292 = 128'b01010001100011000100000001011101110111101001111000011101011111110110010010000000100100000000111001101101000110011010010010110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4292[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4292, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111000010110000110001110000011001001100111110001101010111111011010001001110001111100100100101110100000011101101110101001101110; 
out4293 = 128'b11010101001110001101010011001111100100001001001010111010100111100000011010000111110111001010101000100011001000101000100000101011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4293[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4293, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110000101100001100011100000110010011001111100011010101111110110100010011100011111001001001011101000000111011011101010011011100; 
out4294 = 128'b00111000010001111001100101111111100110010010101110101001100100100110010011010000100010101100100011101011111000101000111000110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4294[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4294, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001011101000000101101011010100000100000101000000100111001111101100111010100011001110111100001001011011101010010001010000011001; 
out4295 = 128'b10011110111011110010100000111000010111010011101010111110101100100111000011011111001011110011110000000011010111000110111111001100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4295[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4295, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010111010000001011010110101000001000001010000001001110011111011001110101000110011101111000010010110111010100100010100000110011; 
out4296 = 128'b00111011111000001100000000110111011111111101110111101010111100001111100111011001101010110100110001100101000010110011101011000011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4296[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4296, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01000100010000001011111110001000110010001110000100010000001100110111110111101000000111011110010110110100110101101110110111000111; 
out4297 = 128'b00111010000011010001100001000101010010010011110111100000001101101101100101000010001011001101001111110011001000110000110100110010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4297[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4297, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001000100000010111111100010001100100011100001000100000011001101111101111010000001110111100101101101001101011011101101110001110; 
out4298 = 128'b00000111001101000001110111001010100100110101001010000110010101010010011111000000111101001010110100010100000011011010011010010001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4298[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4298, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010001000000101111111000100011001000111000010001000000110011011111011110100000011101111001011011010011010110111011011100011100; 
out4299 = 128'b10111111011111011111000101000101000011100111101110010101100010010111100101100111000111000011000011001000110011100000001110001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4299[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4299, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01001000110001000010100010011110110011101010100100001101010100111010100000100100000111011100000101111100110001011101001110011001; 
out4300 = 128'b00100010001101010100110111000101110110111001010001111000111000000010110001110100100101101011001010101100111111111001110110101101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4300[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4300, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111011010010011000010111100101000101001111001110010110011011110001011100101100110010010110111000100011111110010001101010010011; 
out4301 = 128'b11100000001011000011011001101101100010100011111010000011101000000100101100100110110101111000101000011001100100010111100001110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4301[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4301, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11110110100100110000101111001010001010011110011100101100110111100010111001011001100100101101110001000111111100100011010100100110; 
out4302 = 128'b00000111111011000010000110010001001100111011100110101100010010001000001100001000001111011110011011010010011101000101101101001011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4302[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4302, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000111111001111100001101001100110110100110111111010101011101000001101111010111110101110101010001010101100101101101011111101101; 
out4303 = 128'b10110110101111101001100101010100110111001110100111110011010000010001010000000000011100001000111101101001110101000100010011011010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4303[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4303, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001111110011111000011010011001101101001101111110101010111010000011011110101111101011101010100010101011001011011010111111011011; 
out4304 = 128'b00111010100100001010110000100101100111010010001100100011101110010011111000100001011101111100101100000111100011001011000111111010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4304[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4304, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110101010111101101100111101011111000000001111011011001000110000010100000111011101011111011110110001100001010011110001000010110; 
out4305 = 128'b00101101111101111011010111001110100110000111011000010111010010100101011111011011101000100101011101101111010110010001100010110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4305[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4305, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000000011111000110011100001111010010011001110000111110111110000001011100010011101011011001011111000010001000010111100110001100; 
out4306 = 128'b11000101111001000000111101111001010010011101100101000100100010011101001111111111001011111000100011100000011100000010110110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4306[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4306, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000000111110001100111000011110100100110011100001111101111100000010111000100111010110110010111110000100010000101111001100011001; 
out4307 = 128'b00110000110001101001100110110101100101001101001001000101001101001111111001111000010110100000001000000111010011011100100100110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4307[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4307, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000001111100011001110000111101001001100111000011111011111000000101110001001110101101100101111100001000100001011110011000110011; 
out4308 = 128'b10011101001000010110101000001101111001100010111011001111001010000011010001110111001111111110010001100010111011000000110000100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4308[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4308, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000011111000110011100001111010010011001110000111110111110000001011100010011101011011001011111000010001000010111100110001100110; 
out4309 = 128'b01110011000101100110110001111100000001010001011001100100001101111101101101101110010101011010110100000101110001110111011100100010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4309[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4309, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000111110001100111000011110100100110011100001111101111100000010111000100111010110110010111110000100010000101111001100011001101; 
out4310 = 128'b11100110110010001011110010000100100111010111000101100000100001111101100101010010011000111101011101011001001011000100111111111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4310[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4310, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100101010011010011010100110001101110100010011001010011110010101010010100010001010000000001010010011110010111011000110000111011; 
out4311 = 128'b10000100100101100010111101101101011110111010100110011001111111110010011000000101110110110011010110110010001101111101000011111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4311[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4311, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100000010110111011111010111011111111011110110100101011010111010000110101000110011100101100010111100110110010011010010111010111; 
out4312 = 128'b11001100110010011010100100110000110000001001110011111111101010101000100101100110010001111111011001111111011111111111101101111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4312[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4312, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00101010011101101010100110101111011100100111101111011010011100100101110111101000000101110110011100010111111000011111011000001111; 
out4313 = 128'b00001101111000010001010100001011111111000110000011111010010000001110101111110001110001010110010101010001100001111000010000101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4313[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4313, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01010100111011010101001101011110111001001111011110110100111001001011101111010000001011101100111000101111110000111110110000011111; 
out4314 = 128'b00011011100010000100100111000100110111011000111001001000111010001110100010100111110111111100011011100010010110110110001000100111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4314[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4314, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11000011000110110111001001100101010000000100111011100101000000010011000011000100101011110111000010000101111101010110010110011110; 
out4315 = 128'b11011111111000101110110011101111000010110100111010111000010110100111111000011110110100110000001011000010011111101001010100101000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4315[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4315, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10000110001101101110010011001010100000001001110111001010000000100110000110001001010111101110000100001011111010101100101100111101; 
out4316 = 128'b00010100111001011001001010000101111001000101000110101010110000001001001010101111111100100010111111100010111011111100110101100101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4316[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4316, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01100110101011000001110101001101100010001001101000011000110011001000010001110110010011110010111011001101101001110010101111011010; 
out4317 = 128'b11010110010111000011111101010100001101001000001010010110010000010000100001010111010110010111000011011010011001101101000001111111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4317[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4317, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11001101010110000011101010011011000100010011010000110001100110010000100011101100100111100101110110011011010011100101011110110100; 
out4318 = 128'b01001110101010111010100000100101010110101000100011001110011110100101010011000000101001100101110011010010111100101011010111100011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4318[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4318, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10011010101100000111010100110110001000100110100001100011001100100001000111011001001111001011101100110110100111001010111101101000; 
out4319 = 128'b10010011100110110010111010011111000111100011111111111111011001000001100101000000111100111110101001110100100010000101110100000111; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4319[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4319, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00110101011000001110101001101100010001001101000011000110011001000010001110110010011110010111011001101101001110010101111011010000; 
out4320 = 128'b01110100110011010001101111010010001101100110001110001101010001100101110110011011100001000000000111001100100100001011101100000000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4320[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4320, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110100110010010110101110001010000011011010111001110110110010100100100000010000010110011010100111011111101100110100010000111000; 
out4321 = 128'b00101100111110100110001010100111001011111101100011111111100001001001011000111101110010110111101110000011010100110011111110001101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4321[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4321, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11101001100100101101011100010100000110110101110011101101100101001001000000100000101100110101001110111111011001101000100001110001; 
out4322 = 128'b10001111001010100110010011011011011001001010001100100111110110100110100111010101001011010110011010101000100010010101000110111001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4322[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4322, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10100111111011001100010110100010001110110001011110101101111000110110100001010001001111110000111010100001011111100101010011011010; 
out4323 = 128'b11101100010001000000000000000011110111010101010011100110010110000100110100100110111111011011101100011011010100110110010000001001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4323[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4323, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111011000100001110000011001110011110111000000100101101000011001001100010110010001001111011010010011101010011111110110110001101; 
out4324 = 128'b11001111101100001011101110110001111111001111001000010110000100000110101111011000110011110000000011011111000100000000101001101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4324[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4324, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000010111010001010101000010110111110101010110000101100110100110111100101110100000101101100000011100101001011001001111100100011; 
out4325 = 128'b01111011000101111110101101100100111110111000110011010111100111110011010001010001001000011000110011111110000011000000110100001110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4325[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4325, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00000101110100010101010000101101111101010101100001011001101001101111001011101000001011011000000111001010010110010011111001000111; 
out4326 = 128'b00101001001000010010001010000001000010001001110011001100010010101110110001010101011111110101111001101011011010001101001110010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4326[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4326, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01111111011010111100001111010001111001110001111011000101100001111010110111000000000000101010101001001011000000010011100010110110; 
out4327 = 128'b11101001111100010001100100000100110100100011000101000000000000001101010011001111010000100110010101101011000000011111110010100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4327[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4327, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b11111110110101111000011110100011110011100011110110001011000011110101101110000000000001010101010010010110000000100111000101101101; 
out4328 = 128'b11001110101100001110111110010001001100010011010001001000000111101111011001100110101101111111110110111010100000111111011011100000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4328[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4328, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10001001011001100110010011001101100100011101010101100000110101001111111100010000010100110000000011110011101101111010011011100010; 
out4329 = 128'b00001001100100000000110111110100101001001001100000100010110000011001000111010011110011011111000100111001100101000011101001011101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4329[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4329, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010010110011001100100110011011001000111010101011000001101010011111111000100000101001100000000111100111011011110100110111000101; 
out4330 = 128'b10110011101100011010110001101001111001001001000101110101011010101010110100100000010111110011010010000001111001001100011101110100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4330[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4330, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00100101100110011001001100110110010001110101010110000011010100111111110001000001010011000000001111001110110111101001101110001011; 
out4331 = 128'b11101100000101110000000011100101101110001100111001011100101000000001110101001001011111111100011100111010111000000100100011011100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4331[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4331, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00111111111110100100110111100110100000110000010101110000011011011011000010010010110000011010111001000010000011100111001100101110; 
out4332 = 128'b10100101111000001111001100100100000101010000010001001010111011111000001110100110111110010110101010101111010010011111010101110101; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4332[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4332, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00001011001111011111000001000111000010111010010010010110000100010010100100110101110110101111010101011011101011111010001001100100; 
out4333 = 128'b01000010110111010001000110100001001100000110111010001101010110000100000100011100010101011111000010011100010011001111001110000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4333[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4333, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010110011110111110000010001110000101110100100100101100001000100101001001101011101101011110101010110111010111110100010011001001; 
out4334 = 128'b10101010101000101111000000011010000101101110010111110101101000010000001111001001100010110100111010110001001000011110010101101010; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4334[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4334, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011000001111101010101010010110001000110011110000101110100011101110110011000111001100100111110010110001000011011100110110101011; 
out4335 = 128'b00110001001001001011101100001000110001001100110000100000110001011111010001110001010000010001101011100101011111100110011000110000; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4335[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4335, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10110000011111010101010100101100010001100111100001011101000111011101100110001110011001001111100101100010000110111001101101010111; 
out4336 = 128'b11110110011011010011010110101111100001101010011100010100000101010001110101001111001110011110100011001010001101111001001110101001; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4336[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4336, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b00010100001100111100000111010010100000010101111011001100111100011111101100001100100100000101101100011011100001000111001010010110; 
out4337 = 128'b11010111100010111001101101000100110001101011111100000000011010001110101100000100000000100100110110000010000000100001110110110011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4337[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4337, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01011100101011101110100000101111000011110001001111101111001010011011111000001001011110010001111111101000101110111010000100010101; 
out4338 = 128'b00101100011110000001100101001100110001110101101000011000101011111110110000010011001110101100100010111011010110010000100110000100; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4338[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4338, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b10111001010111011101000001011110000111100010011111011110010100110111110000010010111100100011111111010001011101110100001000101010; 
out4339 = 128'b10010111010110010010011100010100100010000111010101000001011100010111111101010010000110100011011101101001001010101011001011010011; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4339[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4339, out, Antena); 
#100; 
@ (negedge clk); 
#2; 
key = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
state = 128'b01110010101110111010000010111100001111000100111110111100101001101111100000100101111001000111111110100010111011101000010001010101; 
out4340 = 128'b00000110110000110001011011000111001100000100100110010000001100011001101001111101101011111110001010101001000000001111011000100110; 
#7.1;
for (i=0;i<128;i=i+1) begin 
if (out[i] != out4340[i]) begin 
bit_err = bit_err + 128'b1; 
end 
end 
$fwrite(f,"%b, %b, %b, %b\n",state, out4340, out, Antena); 
$display("%d", bit_err); 
$fclose(f); 
$finish; 
end 
always #5 clk = ~clk; 
endmodule 
